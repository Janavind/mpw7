VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.490 748.240 426.810 748.300 ;
        RECT 447.190 748.240 447.510 748.300 ;
        RECT 426.490 748.100 447.510 748.240 ;
        RECT 426.490 748.040 426.810 748.100 ;
        RECT 447.190 748.040 447.510 748.100 ;
        RECT 458.230 748.240 458.550 748.300 ;
        RECT 458.230 748.100 496.870 748.240 ;
        RECT 458.230 748.040 458.550 748.100 ;
        RECT 447.190 747.220 447.510 747.280 ;
        RECT 458.230 747.220 458.550 747.280 ;
        RECT 447.190 747.080 458.550 747.220 ;
        RECT 496.730 747.220 496.870 748.100 ;
        RECT 517.430 747.420 614.170 747.560 ;
        RECT 517.430 747.220 517.570 747.420 ;
        RECT 496.730 747.080 517.570 747.220 ;
        RECT 614.030 747.220 614.170 747.420 ;
        RECT 2901.290 747.220 2901.610 747.280 ;
        RECT 614.030 747.080 2901.610 747.220 ;
        RECT 447.190 747.020 447.510 747.080 ;
        RECT 458.230 747.020 458.550 747.080 ;
        RECT 2901.290 747.020 2901.610 747.080 ;
      LAYER via ;
        RECT 426.520 748.040 426.780 748.300 ;
        RECT 447.220 748.040 447.480 748.300 ;
        RECT 458.260 748.040 458.520 748.300 ;
        RECT 447.220 747.020 447.480 747.280 ;
        RECT 458.260 747.020 458.520 747.280 ;
        RECT 2901.320 747.020 2901.580 747.280 ;
      LAYER met2 ;
        RECT 425.850 748.410 426.130 750.000 ;
        RECT 425.850 748.330 426.720 748.410 ;
        RECT 425.850 748.270 426.780 748.330 ;
        RECT 425.850 746.000 426.130 748.270 ;
        RECT 426.520 748.010 426.780 748.270 ;
        RECT 447.220 748.010 447.480 748.330 ;
        RECT 458.260 748.010 458.520 748.330 ;
        RECT 447.280 747.310 447.420 748.010 ;
        RECT 458.320 747.310 458.460 748.010 ;
        RECT 447.220 746.990 447.480 747.310 ;
        RECT 458.260 746.990 458.520 747.310 ;
        RECT 2901.320 746.990 2901.580 747.310 ;
        RECT 2901.380 39.285 2901.520 746.990 ;
        RECT 2901.310 38.915 2901.590 39.285 ;
      LAYER via2 ;
        RECT 2901.310 38.960 2901.590 39.240 ;
      LAYER met3 ;
        RECT 2901.285 39.250 2901.615 39.265 ;
        RECT 2917.600 39.250 2924.800 39.700 ;
        RECT 2901.285 38.950 2924.800 39.250 ;
        RECT 2901.285 38.935 2901.615 38.950 ;
        RECT 2917.600 38.500 2924.800 38.950 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.550 2380.580 477.870 2380.640 ;
        RECT 2900.830 2380.580 2901.150 2380.640 ;
        RECT 477.550 2380.440 2901.150 2380.580 ;
        RECT 477.550 2380.380 477.870 2380.440 ;
        RECT 2900.830 2380.380 2901.150 2380.440 ;
        RECT 477.550 766.600 477.870 766.660 ;
        RECT 480.310 766.600 480.630 766.660 ;
        RECT 477.550 766.460 480.630 766.600 ;
        RECT 477.550 766.400 477.870 766.460 ;
        RECT 480.310 766.400 480.630 766.460 ;
      LAYER via ;
        RECT 477.580 2380.380 477.840 2380.640 ;
        RECT 2900.860 2380.380 2901.120 2380.640 ;
        RECT 477.580 766.400 477.840 766.660 ;
        RECT 480.340 766.400 480.600 766.660 ;
      LAYER met2 ;
        RECT 2900.850 2384.915 2901.130 2385.285 ;
        RECT 2900.920 2380.670 2901.060 2384.915 ;
        RECT 477.580 2380.350 477.840 2380.670 ;
        RECT 2900.860 2380.350 2901.120 2380.670 ;
        RECT 477.640 766.690 477.780 2380.350 ;
        RECT 477.580 766.370 477.840 766.690 ;
        RECT 480.340 766.370 480.600 766.690 ;
        RECT 480.400 749.770 480.540 766.370 ;
        RECT 481.050 749.770 481.330 750.000 ;
        RECT 480.400 749.630 481.330 749.770 ;
        RECT 481.050 746.000 481.330 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2384.960 2901.130 2385.240 ;
      LAYER met3 ;
        RECT 2900.825 2385.250 2901.155 2385.265 ;
        RECT 2917.600 2385.250 2924.800 2385.700 ;
        RECT 2900.825 2384.950 2924.800 2385.250 ;
        RECT 2900.825 2384.935 2901.155 2384.950 ;
        RECT 2917.600 2384.500 2924.800 2384.950 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 485.830 2615.180 486.150 2615.240 ;
        RECT 2900.830 2615.180 2901.150 2615.240 ;
        RECT 485.830 2615.040 2901.150 2615.180 ;
        RECT 485.830 2614.980 486.150 2615.040 ;
        RECT 2900.830 2614.980 2901.150 2615.040 ;
      LAYER via ;
        RECT 485.860 2614.980 486.120 2615.240 ;
        RECT 2900.860 2614.980 2901.120 2615.240 ;
      LAYER met2 ;
        RECT 2900.850 2619.515 2901.130 2619.885 ;
        RECT 2900.920 2615.270 2901.060 2619.515 ;
        RECT 485.860 2614.950 486.120 2615.270 ;
        RECT 2900.860 2614.950 2901.120 2615.270 ;
        RECT 485.920 749.770 486.060 2614.950 ;
        RECT 486.570 749.770 486.850 750.000 ;
        RECT 485.920 749.630 486.850 749.770 ;
        RECT 486.570 746.000 486.850 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2619.560 2901.130 2619.840 ;
      LAYER met3 ;
        RECT 2900.825 2619.850 2901.155 2619.865 ;
        RECT 2917.600 2619.850 2924.800 2620.300 ;
        RECT 2900.825 2619.550 2924.800 2619.850 ;
        RECT 2900.825 2619.535 2901.155 2619.550 ;
        RECT 2917.600 2619.100 2924.800 2619.550 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.810 2849.780 492.130 2849.840 ;
        RECT 2900.830 2849.780 2901.150 2849.840 ;
        RECT 491.810 2849.640 2901.150 2849.780 ;
        RECT 491.810 2849.580 492.130 2849.640 ;
        RECT 2900.830 2849.580 2901.150 2849.640 ;
      LAYER via ;
        RECT 491.840 2849.580 492.100 2849.840 ;
        RECT 2900.860 2849.580 2901.120 2849.840 ;
      LAYER met2 ;
        RECT 2900.850 2854.115 2901.130 2854.485 ;
        RECT 2900.920 2849.870 2901.060 2854.115 ;
        RECT 491.840 2849.550 492.100 2849.870 ;
        RECT 2900.860 2849.550 2901.120 2849.870 ;
        RECT 491.900 751.130 492.040 2849.550 ;
        RECT 491.900 750.990 492.270 751.130 ;
        RECT 492.130 750.000 492.270 750.990 ;
        RECT 492.090 746.000 492.370 750.000 ;
      LAYER via2 ;
        RECT 2900.850 2854.160 2901.130 2854.440 ;
      LAYER met3 ;
        RECT 2900.825 2854.450 2901.155 2854.465 ;
        RECT 2917.600 2854.450 2924.800 2854.900 ;
        RECT 2900.825 2854.150 2924.800 2854.450 ;
        RECT 2900.825 2854.135 2901.155 2854.150 ;
        RECT 2917.600 2853.700 2924.800 2854.150 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 3084.380 497.650 3084.440 ;
        RECT 2900.830 3084.380 2901.150 3084.440 ;
        RECT 497.330 3084.240 2901.150 3084.380 ;
        RECT 497.330 3084.180 497.650 3084.240 ;
        RECT 2900.830 3084.180 2901.150 3084.240 ;
      LAYER via ;
        RECT 497.360 3084.180 497.620 3084.440 ;
        RECT 2900.860 3084.180 2901.120 3084.440 ;
      LAYER met2 ;
        RECT 2900.850 3088.715 2901.130 3089.085 ;
        RECT 2900.920 3084.470 2901.060 3088.715 ;
        RECT 497.360 3084.150 497.620 3084.470 ;
        RECT 2900.860 3084.150 2901.120 3084.470 ;
        RECT 497.420 751.130 497.560 3084.150 ;
        RECT 497.420 750.990 497.790 751.130 ;
        RECT 497.650 750.000 497.790 750.990 ;
        RECT 497.610 746.000 497.890 750.000 ;
      LAYER via2 ;
        RECT 2900.850 3088.760 2901.130 3089.040 ;
      LAYER met3 ;
        RECT 2900.825 3089.050 2901.155 3089.065 ;
        RECT 2917.600 3089.050 2924.800 3089.500 ;
        RECT 2900.825 3088.750 2924.800 3089.050 ;
        RECT 2900.825 3088.735 2901.155 3088.750 ;
        RECT 2917.600 3088.300 2924.800 3088.750 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 501.010 3318.980 501.330 3319.040 ;
        RECT 2900.830 3318.980 2901.150 3319.040 ;
        RECT 501.010 3318.840 2901.150 3318.980 ;
        RECT 501.010 3318.780 501.330 3318.840 ;
        RECT 2900.830 3318.780 2901.150 3318.840 ;
      LAYER via ;
        RECT 501.040 3318.780 501.300 3319.040 ;
        RECT 2900.860 3318.780 2901.120 3319.040 ;
      LAYER met2 ;
        RECT 2900.850 3323.315 2901.130 3323.685 ;
        RECT 2900.920 3319.070 2901.060 3323.315 ;
        RECT 501.040 3318.750 501.300 3319.070 ;
        RECT 2900.860 3318.750 2901.120 3319.070 ;
        RECT 501.100 855.670 501.240 3318.750 ;
        RECT 501.100 855.530 502.620 855.670 ;
        RECT 502.480 749.770 502.620 855.530 ;
        RECT 503.130 749.770 503.410 750.000 ;
        RECT 502.480 749.630 503.410 749.770 ;
        RECT 503.130 746.000 503.410 749.630 ;
      LAYER via2 ;
        RECT 2900.850 3323.360 2901.130 3323.640 ;
      LAYER met3 ;
        RECT 2900.825 3323.650 2901.155 3323.665 ;
        RECT 2917.600 3323.650 2924.800 3324.100 ;
        RECT 2900.825 3323.350 2924.800 3323.650 ;
        RECT 2900.825 3323.335 2901.155 3323.350 ;
        RECT 2917.600 3322.900 2924.800 3323.350 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.830 769.320 509.150 769.380 ;
        RECT 2863.570 769.320 2863.890 769.380 ;
        RECT 508.830 769.180 2863.890 769.320 ;
        RECT 508.830 769.120 509.150 769.180 ;
        RECT 2863.570 769.120 2863.890 769.180 ;
      LAYER via ;
        RECT 508.860 769.120 509.120 769.380 ;
        RECT 2863.600 769.120 2863.860 769.380 ;
      LAYER met2 ;
        RECT 2864.830 3517.600 2865.390 3524.800 ;
        RECT 2865.040 3512.170 2865.180 3517.600 ;
        RECT 2863.660 3512.030 2865.180 3512.170 ;
        RECT 2863.660 769.410 2863.800 3512.030 ;
        RECT 508.860 769.090 509.120 769.410 ;
        RECT 2863.600 769.090 2863.860 769.410 ;
        RECT 508.920 750.000 509.060 769.090 ;
        RECT 508.650 749.630 509.060 750.000 ;
        RECT 508.650 746.000 508.930 749.630 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.350 769.660 514.670 769.720 ;
        RECT 2539.270 769.660 2539.590 769.720 ;
        RECT 514.350 769.520 2539.590 769.660 ;
        RECT 514.350 769.460 514.670 769.520 ;
        RECT 2539.270 769.460 2539.590 769.520 ;
      LAYER via ;
        RECT 514.380 769.460 514.640 769.720 ;
        RECT 2539.300 769.460 2539.560 769.720 ;
      LAYER met2 ;
        RECT 2540.530 3517.600 2541.090 3524.800 ;
        RECT 2540.740 3512.170 2540.880 3517.600 ;
        RECT 2539.360 3512.030 2540.880 3512.170 ;
        RECT 2539.360 769.750 2539.500 3512.030 ;
        RECT 514.380 769.430 514.640 769.750 ;
        RECT 2539.300 769.430 2539.560 769.750 ;
        RECT 514.440 750.000 514.580 769.430 ;
        RECT 514.170 749.630 514.580 750.000 ;
        RECT 514.170 746.000 514.450 749.630 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.870 770.000 520.190 770.060 ;
        RECT 2214.970 770.000 2215.290 770.060 ;
        RECT 519.870 769.860 2215.290 770.000 ;
        RECT 519.870 769.800 520.190 769.860 ;
        RECT 2214.970 769.800 2215.290 769.860 ;
      LAYER via ;
        RECT 519.900 769.800 520.160 770.060 ;
        RECT 2215.000 769.800 2215.260 770.060 ;
      LAYER met2 ;
        RECT 2216.230 3517.600 2216.790 3524.800 ;
        RECT 2216.440 3512.170 2216.580 3517.600 ;
        RECT 2215.060 3512.030 2216.580 3512.170 ;
        RECT 2215.060 770.090 2215.200 3512.030 ;
        RECT 519.900 769.770 520.160 770.090 ;
        RECT 2215.000 769.770 2215.260 770.090 ;
        RECT 519.960 750.000 520.100 769.770 ;
        RECT 519.690 749.630 520.100 750.000 ;
        RECT 519.690 746.000 519.970 749.630 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 770.340 525.250 770.400 ;
        RECT 1890.670 770.340 1890.990 770.400 ;
        RECT 524.930 770.200 1890.990 770.340 ;
        RECT 524.930 770.140 525.250 770.200 ;
        RECT 1890.670 770.140 1890.990 770.200 ;
      LAYER via ;
        RECT 524.960 770.140 525.220 770.400 ;
        RECT 1890.700 770.140 1890.960 770.400 ;
      LAYER met2 ;
        RECT 1891.930 3517.600 1892.490 3524.800 ;
        RECT 1892.140 3512.170 1892.280 3517.600 ;
        RECT 1890.760 3512.030 1892.280 3512.170 ;
        RECT 1890.760 770.430 1890.900 3512.030 ;
        RECT 524.960 770.110 525.220 770.430 ;
        RECT 1890.700 770.110 1890.960 770.430 ;
        RECT 525.020 751.130 525.160 770.110 ;
        RECT 525.020 750.990 525.390 751.130 ;
        RECT 525.250 750.000 525.390 750.990 ;
        RECT 525.210 746.000 525.490 750.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 530.910 770.680 531.230 770.740 ;
        RECT 1566.370 770.680 1566.690 770.740 ;
        RECT 530.910 770.540 1566.690 770.680 ;
        RECT 530.910 770.480 531.230 770.540 ;
        RECT 1566.370 770.480 1566.690 770.540 ;
      LAYER via ;
        RECT 530.940 770.480 531.200 770.740 ;
        RECT 1566.400 770.480 1566.660 770.740 ;
      LAYER met2 ;
        RECT 1567.630 3517.600 1568.190 3524.800 ;
        RECT 1567.840 3512.170 1567.980 3517.600 ;
        RECT 1566.460 3512.030 1567.980 3512.170 ;
        RECT 1566.460 770.770 1566.600 3512.030 ;
        RECT 530.940 770.450 531.200 770.770 ;
        RECT 1566.400 770.450 1566.660 770.770 ;
        RECT 531.000 750.000 531.140 770.450 ;
        RECT 530.730 749.630 531.140 750.000 ;
        RECT 530.730 746.000 531.010 749.630 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.010 747.020 432.330 747.280 ;
        RECT 432.100 746.880 432.240 747.020 ;
        RECT 431.640 746.740 432.240 746.880 ;
        RECT 431.640 745.860 431.780 746.740 ;
        RECT 2902.210 745.860 2902.530 745.920 ;
        RECT 431.640 745.720 2902.530 745.860 ;
        RECT 2902.210 745.660 2902.530 745.720 ;
      LAYER via ;
        RECT 432.040 747.020 432.300 747.280 ;
        RECT 2902.240 745.660 2902.500 745.920 ;
      LAYER met2 ;
        RECT 431.370 747.050 431.650 750.000 ;
        RECT 432.040 747.050 432.300 747.310 ;
        RECT 431.370 746.990 432.300 747.050 ;
        RECT 431.370 746.910 432.240 746.990 ;
        RECT 431.370 746.000 431.650 746.910 ;
        RECT 2902.240 745.630 2902.500 745.950 ;
        RECT 2902.300 273.885 2902.440 745.630 ;
        RECT 2902.230 273.515 2902.510 273.885 ;
      LAYER via2 ;
        RECT 2902.230 273.560 2902.510 273.840 ;
      LAYER met3 ;
        RECT 2902.205 273.850 2902.535 273.865 ;
        RECT 2917.600 273.850 2924.800 274.300 ;
        RECT 2902.205 273.550 2924.800 273.850 ;
        RECT 2902.205 273.535 2902.535 273.550 ;
        RECT 2917.600 273.100 2924.800 273.550 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.510 777.140 535.830 777.200 ;
        RECT 1242.070 777.140 1242.390 777.200 ;
        RECT 535.510 777.000 1242.390 777.140 ;
        RECT 535.510 776.940 535.830 777.000 ;
        RECT 1242.070 776.940 1242.390 777.000 ;
      LAYER via ;
        RECT 535.540 776.940 535.800 777.200 ;
        RECT 1242.100 776.940 1242.360 777.200 ;
      LAYER met2 ;
        RECT 1243.330 3517.600 1243.890 3524.800 ;
        RECT 1243.540 3512.170 1243.680 3517.600 ;
        RECT 1242.160 3512.030 1243.680 3512.170 ;
        RECT 1242.160 777.230 1242.300 3512.030 ;
        RECT 535.540 776.910 535.800 777.230 ;
        RECT 1242.100 776.910 1242.360 777.230 ;
        RECT 535.600 749.770 535.740 776.910 ;
        RECT 536.250 749.770 536.530 750.000 ;
        RECT 535.600 749.630 536.530 749.770 ;
        RECT 536.250 746.000 536.530 749.630 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.030 778.160 541.350 778.220 ;
        RECT 917.770 778.160 918.090 778.220 ;
        RECT 541.030 778.020 918.090 778.160 ;
        RECT 541.030 777.960 541.350 778.020 ;
        RECT 917.770 777.960 918.090 778.020 ;
      LAYER via ;
        RECT 541.060 777.960 541.320 778.220 ;
        RECT 917.800 777.960 918.060 778.220 ;
      LAYER met2 ;
        RECT 919.030 3517.600 919.590 3524.800 ;
        RECT 919.240 3512.170 919.380 3517.600 ;
        RECT 917.860 3512.030 919.380 3512.170 ;
        RECT 917.860 778.250 918.000 3512.030 ;
        RECT 541.060 777.930 541.320 778.250 ;
        RECT 917.800 777.930 918.060 778.250 ;
        RECT 541.120 749.770 541.260 777.930 ;
        RECT 541.770 749.770 542.050 750.000 ;
        RECT 541.120 749.630 542.050 749.770 ;
        RECT 541.770 746.000 542.050 749.630 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 547.930 771.360 548.250 771.420 ;
        RECT 593.930 771.360 594.250 771.420 ;
        RECT 547.930 771.220 594.250 771.360 ;
        RECT 547.930 771.160 548.250 771.220 ;
        RECT 593.930 771.160 594.250 771.220 ;
      LAYER via ;
        RECT 547.960 771.160 548.220 771.420 ;
        RECT 593.960 771.160 594.220 771.420 ;
      LAYER met2 ;
        RECT 594.730 3517.600 595.290 3524.800 ;
        RECT 594.940 3512.170 595.080 3517.600 ;
        RECT 593.560 3512.030 595.080 3512.170 ;
        RECT 593.560 855.670 593.700 3512.030 ;
        RECT 593.560 855.530 594.160 855.670 ;
        RECT 594.020 771.450 594.160 855.530 ;
        RECT 547.960 771.130 548.220 771.450 ;
        RECT 593.960 771.130 594.220 771.450 ;
        RECT 547.290 749.770 547.570 750.000 ;
        RECT 548.020 749.770 548.160 771.130 ;
        RECT 547.290 749.630 548.160 749.770 ;
        RECT 547.290 746.000 547.570 749.630 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.170 771.020 269.490 771.080 ;
        RECT 552.070 771.020 552.390 771.080 ;
        RECT 269.170 770.880 552.390 771.020 ;
        RECT 269.170 770.820 269.490 770.880 ;
        RECT 552.070 770.820 552.390 770.880 ;
      LAYER via ;
        RECT 269.200 770.820 269.460 771.080 ;
        RECT 552.100 770.820 552.360 771.080 ;
      LAYER met2 ;
        RECT 270.430 3517.600 270.990 3524.800 ;
        RECT 270.640 3512.170 270.780 3517.600 ;
        RECT 269.260 3512.030 270.780 3512.170 ;
        RECT 269.260 771.110 269.400 3512.030 ;
        RECT 269.200 770.790 269.460 771.110 ;
        RECT 552.100 770.790 552.360 771.110 ;
        RECT 552.160 749.770 552.300 770.790 ;
        RECT 552.810 749.770 553.090 750.000 ;
        RECT 552.160 749.630 553.090 749.770 ;
        RECT 552.810 746.000 553.090 749.630 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3470.960 17.410 3471.020 ;
        RECT 556.210 3470.960 556.530 3471.020 ;
        RECT 17.090 3470.820 556.530 3470.960 ;
        RECT 17.090 3470.760 17.410 3470.820 ;
        RECT 556.210 3470.760 556.530 3470.820 ;
      LAYER via ;
        RECT 17.120 3470.760 17.380 3471.020 ;
        RECT 556.240 3470.760 556.500 3471.020 ;
      LAYER met2 ;
        RECT 17.110 3474.275 17.390 3474.645 ;
        RECT 17.180 3471.050 17.320 3474.275 ;
        RECT 17.120 3470.730 17.380 3471.050 ;
        RECT 556.240 3470.730 556.500 3471.050 ;
        RECT 556.300 855.670 556.440 3470.730 ;
        RECT 556.300 855.530 557.820 855.670 ;
        RECT 557.680 749.770 557.820 855.530 ;
        RECT 558.330 749.770 558.610 750.000 ;
        RECT 557.680 749.630 558.610 749.770 ;
        RECT 558.330 746.000 558.610 749.630 ;
      LAYER via2 ;
        RECT 17.110 3474.320 17.390 3474.600 ;
      LAYER met3 ;
        RECT -4.800 3474.610 2.400 3475.060 ;
        RECT 17.085 3474.610 17.415 3474.625 ;
        RECT -4.800 3474.310 17.415 3474.610 ;
        RECT -4.800 3473.860 2.400 3474.310 ;
        RECT 17.085 3474.295 17.415 3474.310 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 3222.420 16.490 3222.480 ;
        RECT 561.730 3222.420 562.050 3222.480 ;
        RECT 16.170 3222.280 562.050 3222.420 ;
        RECT 16.170 3222.220 16.490 3222.280 ;
        RECT 561.730 3222.220 562.050 3222.280 ;
        RECT 561.730 749.260 562.050 749.320 ;
        RECT 563.110 749.260 563.430 749.320 ;
        RECT 561.730 749.120 563.430 749.260 ;
        RECT 561.730 749.060 562.050 749.120 ;
        RECT 563.110 749.060 563.430 749.120 ;
      LAYER via ;
        RECT 16.200 3222.220 16.460 3222.480 ;
        RECT 561.760 3222.220 562.020 3222.480 ;
        RECT 561.760 749.060 562.020 749.320 ;
        RECT 563.140 749.060 563.400 749.320 ;
      LAYER met2 ;
        RECT 16.190 3223.355 16.470 3223.725 ;
        RECT 16.260 3222.510 16.400 3223.355 ;
        RECT 16.200 3222.190 16.460 3222.510 ;
        RECT 561.760 3222.190 562.020 3222.510 ;
        RECT 561.820 749.350 561.960 3222.190 ;
        RECT 561.760 749.030 562.020 749.350 ;
        RECT 563.140 749.090 563.400 749.350 ;
        RECT 563.850 749.090 564.130 750.000 ;
        RECT 563.140 749.030 564.130 749.090 ;
        RECT 563.200 748.950 564.130 749.030 ;
        RECT 563.850 746.000 564.130 748.950 ;
      LAYER via2 ;
        RECT 16.190 3223.400 16.470 3223.680 ;
      LAYER met3 ;
        RECT -4.800 3223.690 2.400 3224.140 ;
        RECT 16.165 3223.690 16.495 3223.705 ;
        RECT -4.800 3223.390 16.495 3223.690 ;
        RECT -4.800 3222.940 2.400 3223.390 ;
        RECT 16.165 3223.375 16.495 3223.390 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 777.820 17.410 777.880 ;
        RECT 568.630 777.820 568.950 777.880 ;
        RECT 17.090 777.680 568.950 777.820 ;
        RECT 17.090 777.620 17.410 777.680 ;
        RECT 568.630 777.620 568.950 777.680 ;
      LAYER via ;
        RECT 17.120 777.620 17.380 777.880 ;
        RECT 568.660 777.620 568.920 777.880 ;
      LAYER met2 ;
        RECT 17.110 2972.435 17.390 2972.805 ;
        RECT 17.180 777.910 17.320 2972.435 ;
        RECT 17.120 777.590 17.380 777.910 ;
        RECT 568.660 777.590 568.920 777.910 ;
        RECT 568.720 749.770 568.860 777.590 ;
        RECT 569.370 749.770 569.650 750.000 ;
        RECT 568.720 749.630 569.650 749.770 ;
        RECT 569.370 746.000 569.650 749.630 ;
      LAYER via2 ;
        RECT 17.110 2972.480 17.390 2972.760 ;
      LAYER met3 ;
        RECT -4.800 2972.770 2.400 2973.220 ;
        RECT 17.085 2972.770 17.415 2972.785 ;
        RECT -4.800 2972.470 17.415 2972.770 ;
        RECT -4.800 2972.020 2.400 2972.470 ;
        RECT 17.085 2972.455 17.415 2972.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 777.480 17.870 777.540 ;
        RECT 574.610 777.480 574.930 777.540 ;
        RECT 17.550 777.340 574.930 777.480 ;
        RECT 17.550 777.280 17.870 777.340 ;
        RECT 574.610 777.280 574.930 777.340 ;
      LAYER via ;
        RECT 17.580 777.280 17.840 777.540 ;
        RECT 574.640 777.280 574.900 777.540 ;
      LAYER met2 ;
        RECT 17.570 2721.515 17.850 2721.885 ;
        RECT 17.640 777.570 17.780 2721.515 ;
        RECT 17.580 777.250 17.840 777.570 ;
        RECT 574.640 777.250 574.900 777.570 ;
        RECT 574.700 751.130 574.840 777.250 ;
        RECT 574.700 750.990 575.070 751.130 ;
        RECT 574.930 750.000 575.070 750.990 ;
        RECT 574.890 746.000 575.170 750.000 ;
      LAYER via2 ;
        RECT 17.570 2721.560 17.850 2721.840 ;
      LAYER met3 ;
        RECT -4.800 2721.850 2.400 2722.300 ;
        RECT 17.545 2721.850 17.875 2721.865 ;
        RECT -4.800 2721.550 17.875 2721.850 ;
        RECT -4.800 2721.100 2.400 2721.550 ;
        RECT 17.545 2721.535 17.875 2721.550 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2470.340 16.950 2470.400 ;
        RECT 582.430 2470.340 582.750 2470.400 ;
        RECT 16.630 2470.200 582.750 2470.340 ;
        RECT 16.630 2470.140 16.950 2470.200 ;
        RECT 582.430 2470.140 582.750 2470.200 ;
      LAYER via ;
        RECT 16.660 2470.140 16.920 2470.400 ;
        RECT 582.460 2470.140 582.720 2470.400 ;
      LAYER met2 ;
        RECT 16.650 2470.595 16.930 2470.965 ;
        RECT 16.720 2470.430 16.860 2470.595 ;
        RECT 16.660 2470.110 16.920 2470.430 ;
        RECT 582.460 2470.110 582.720 2470.430 ;
        RECT 582.520 807.370 582.660 2470.110 ;
        RECT 581.140 807.230 582.660 807.370 ;
        RECT 580.410 749.770 580.690 750.000 ;
        RECT 581.140 749.770 581.280 807.230 ;
        RECT 580.410 749.630 581.280 749.770 ;
        RECT 580.410 746.000 580.690 749.630 ;
      LAYER via2 ;
        RECT 16.650 2470.640 16.930 2470.920 ;
      LAYER met3 ;
        RECT -4.800 2470.930 2.400 2471.380 ;
        RECT 16.625 2470.930 16.955 2470.945 ;
        RECT -4.800 2470.630 16.955 2470.930 ;
        RECT -4.800 2470.180 2.400 2470.630 ;
        RECT 16.625 2470.615 16.955 2470.630 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2215.000 16.950 2215.060 ;
        RECT 585.190 2215.000 585.510 2215.060 ;
        RECT 16.630 2214.860 585.510 2215.000 ;
        RECT 16.630 2214.800 16.950 2214.860 ;
        RECT 585.190 2214.800 585.510 2214.860 ;
      LAYER via ;
        RECT 16.660 2214.800 16.920 2215.060 ;
        RECT 585.220 2214.800 585.480 2215.060 ;
      LAYER met2 ;
        RECT 16.650 2219.675 16.930 2220.045 ;
        RECT 16.720 2215.090 16.860 2219.675 ;
        RECT 16.660 2214.770 16.920 2215.090 ;
        RECT 585.220 2214.770 585.480 2215.090 ;
        RECT 585.280 749.770 585.420 2214.770 ;
        RECT 585.930 749.770 586.210 750.000 ;
        RECT 585.280 749.630 586.210 749.770 ;
        RECT 585.930 746.000 586.210 749.630 ;
      LAYER via2 ;
        RECT 16.650 2219.720 16.930 2220.000 ;
      LAYER met3 ;
        RECT -4.800 2220.010 2.400 2220.460 ;
        RECT 16.625 2220.010 16.955 2220.025 ;
        RECT -4.800 2219.710 16.955 2220.010 ;
        RECT -4.800 2219.260 2.400 2219.710 ;
        RECT 16.625 2219.695 16.955 2219.710 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.650 747.020 470.970 747.280 ;
        RECT 470.740 746.540 470.880 747.020 ;
        RECT 2903.130 746.540 2903.450 746.600 ;
        RECT 470.740 746.400 2903.450 746.540 ;
        RECT 2903.130 746.340 2903.450 746.400 ;
      LAYER via ;
        RECT 470.680 747.020 470.940 747.280 ;
        RECT 2903.160 746.340 2903.420 746.600 ;
      LAYER met2 ;
        RECT 436.890 747.730 437.170 750.000 ;
        RECT 437.550 747.730 437.830 747.845 ;
        RECT 436.890 747.590 437.830 747.730 ;
        RECT 436.890 746.000 437.170 747.590 ;
        RECT 437.550 747.475 437.830 747.590 ;
        RECT 470.670 747.475 470.950 747.845 ;
        RECT 470.740 747.310 470.880 747.475 ;
        RECT 470.680 746.990 470.940 747.310 ;
        RECT 2903.160 746.310 2903.420 746.630 ;
        RECT 2903.220 508.485 2903.360 746.310 ;
        RECT 2903.150 508.115 2903.430 508.485 ;
      LAYER via2 ;
        RECT 437.550 747.520 437.830 747.800 ;
        RECT 470.670 747.520 470.950 747.800 ;
        RECT 2903.150 508.160 2903.430 508.440 ;
      LAYER met3 ;
        RECT 437.525 747.810 437.855 747.825 ;
        RECT 470.645 747.810 470.975 747.825 ;
        RECT 437.525 747.510 470.975 747.810 ;
        RECT 437.525 747.495 437.855 747.510 ;
        RECT 470.645 747.495 470.975 747.510 ;
        RECT 2903.125 508.450 2903.455 508.465 ;
        RECT 2917.600 508.450 2924.800 508.900 ;
        RECT 2903.125 508.150 2924.800 508.450 ;
        RECT 2903.125 508.135 2903.455 508.150 ;
        RECT 2917.600 507.700 2924.800 508.150 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1966.800 18.330 1966.860 ;
        RECT 589.330 1966.800 589.650 1966.860 ;
        RECT 18.010 1966.660 589.650 1966.800 ;
        RECT 18.010 1966.600 18.330 1966.660 ;
        RECT 589.330 1966.600 589.650 1966.660 ;
      LAYER via ;
        RECT 18.040 1966.600 18.300 1966.860 ;
        RECT 589.360 1966.600 589.620 1966.860 ;
      LAYER met2 ;
        RECT 18.030 1968.755 18.310 1969.125 ;
        RECT 18.100 1966.890 18.240 1968.755 ;
        RECT 18.040 1966.570 18.300 1966.890 ;
        RECT 589.360 1966.570 589.620 1966.890 ;
        RECT 589.420 759.070 589.560 1966.570 ;
        RECT 589.420 758.930 590.940 759.070 ;
        RECT 590.800 749.770 590.940 758.930 ;
        RECT 591.450 749.770 591.730 750.000 ;
        RECT 590.800 749.630 591.730 749.770 ;
        RECT 591.450 746.000 591.730 749.630 ;
      LAYER via2 ;
        RECT 18.030 1968.800 18.310 1969.080 ;
      LAYER met3 ;
        RECT -4.800 1969.090 2.400 1969.540 ;
        RECT 18.005 1969.090 18.335 1969.105 ;
        RECT -4.800 1968.790 18.335 1969.090 ;
        RECT -4.800 1968.340 2.400 1968.790 ;
        RECT 18.005 1968.775 18.335 1968.790 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1711.460 16.950 1711.520 ;
        RECT 596.690 1711.460 597.010 1711.520 ;
        RECT 16.630 1711.320 597.010 1711.460 ;
        RECT 16.630 1711.260 16.950 1711.320 ;
        RECT 596.690 1711.260 597.010 1711.320 ;
      LAYER via ;
        RECT 16.660 1711.260 16.920 1711.520 ;
        RECT 596.720 1711.260 596.980 1711.520 ;
      LAYER met2 ;
        RECT 16.650 1717.835 16.930 1718.205 ;
        RECT 16.720 1711.550 16.860 1717.835 ;
        RECT 16.660 1711.230 16.920 1711.550 ;
        RECT 596.720 1711.230 596.980 1711.550 ;
        RECT 596.780 751.130 596.920 1711.230 ;
        RECT 596.780 750.990 597.150 751.130 ;
        RECT 597.010 750.000 597.150 750.990 ;
        RECT 596.970 746.000 597.250 750.000 ;
      LAYER via2 ;
        RECT 16.650 1717.880 16.930 1718.160 ;
      LAYER met3 ;
        RECT -4.800 1718.170 2.400 1718.620 ;
        RECT 16.625 1718.170 16.955 1718.185 ;
        RECT -4.800 1717.870 16.955 1718.170 ;
        RECT -4.800 1717.420 2.400 1717.870 ;
        RECT 16.625 1717.855 16.955 1717.870 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1462.920 16.950 1462.980 ;
        RECT 603.130 1462.920 603.450 1462.980 ;
        RECT 16.630 1462.780 603.450 1462.920 ;
        RECT 16.630 1462.720 16.950 1462.780 ;
        RECT 603.130 1462.720 603.450 1462.780 ;
        RECT 601.750 782.920 602.070 782.980 ;
        RECT 603.130 782.920 603.450 782.980 ;
        RECT 601.750 782.780 603.450 782.920 ;
        RECT 601.750 782.720 602.070 782.780 ;
        RECT 603.130 782.720 603.450 782.780 ;
      LAYER via ;
        RECT 16.660 1462.720 16.920 1462.980 ;
        RECT 603.160 1462.720 603.420 1462.980 ;
        RECT 601.780 782.720 602.040 782.980 ;
        RECT 603.160 782.720 603.420 782.980 ;
      LAYER met2 ;
        RECT 16.650 1466.915 16.930 1467.285 ;
        RECT 16.720 1463.010 16.860 1466.915 ;
        RECT 16.660 1462.690 16.920 1463.010 ;
        RECT 603.160 1462.690 603.420 1463.010 ;
        RECT 603.220 783.010 603.360 1462.690 ;
        RECT 601.780 782.690 602.040 783.010 ;
        RECT 603.160 782.690 603.420 783.010 ;
        RECT 601.110 749.770 601.390 750.000 ;
        RECT 601.840 749.770 601.980 782.690 ;
        RECT 601.110 749.630 601.980 749.770 ;
        RECT 601.110 746.000 601.390 749.630 ;
      LAYER via2 ;
        RECT 16.650 1466.960 16.930 1467.240 ;
      LAYER met3 ;
        RECT -4.800 1467.250 2.400 1467.700 ;
        RECT 16.625 1467.250 16.955 1467.265 ;
        RECT -4.800 1466.950 16.955 1467.250 ;
        RECT -4.800 1466.500 2.400 1466.950 ;
        RECT 16.625 1466.935 16.955 1466.950 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1214.720 16.950 1214.780 ;
        RECT 601.750 1214.720 602.070 1214.780 ;
        RECT 16.630 1214.580 602.070 1214.720 ;
        RECT 16.630 1214.520 16.950 1214.580 ;
        RECT 601.750 1214.520 602.070 1214.580 ;
        RECT 601.750 784.280 602.070 784.340 ;
        RECT 604.510 784.280 604.830 784.340 ;
        RECT 601.750 784.140 604.830 784.280 ;
        RECT 601.750 784.080 602.070 784.140 ;
        RECT 604.510 784.080 604.830 784.140 ;
      LAYER via ;
        RECT 16.660 1214.520 16.920 1214.780 ;
        RECT 601.780 1214.520 602.040 1214.780 ;
        RECT 601.780 784.080 602.040 784.340 ;
        RECT 604.540 784.080 604.800 784.340 ;
      LAYER met2 ;
        RECT 16.650 1215.995 16.930 1216.365 ;
        RECT 16.720 1214.810 16.860 1215.995 ;
        RECT 16.660 1214.490 16.920 1214.810 ;
        RECT 601.780 1214.490 602.040 1214.810 ;
        RECT 601.840 784.370 601.980 1214.490 ;
        RECT 601.780 784.050 602.040 784.370 ;
        RECT 604.540 784.050 604.800 784.370 ;
        RECT 604.600 749.770 604.740 784.050 ;
        RECT 605.250 749.770 605.530 750.000 ;
        RECT 604.600 749.630 605.530 749.770 ;
        RECT 605.250 746.000 605.530 749.630 ;
      LAYER via2 ;
        RECT 16.650 1216.040 16.930 1216.320 ;
      LAYER met3 ;
        RECT -4.800 1216.330 2.400 1216.780 ;
        RECT 16.625 1216.330 16.955 1216.345 ;
        RECT -4.800 1216.030 16.955 1216.330 ;
        RECT -4.800 1215.580 2.400 1216.030 ;
        RECT 16.625 1216.015 16.955 1216.030 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 959.380 16.950 959.440 ;
        RECT 608.650 959.380 608.970 959.440 ;
        RECT 16.630 959.240 608.970 959.380 ;
        RECT 16.630 959.180 16.950 959.240 ;
        RECT 608.650 959.180 608.970 959.240 ;
      LAYER via ;
        RECT 16.660 959.180 16.920 959.440 ;
        RECT 608.680 959.180 608.940 959.440 ;
      LAYER met2 ;
        RECT 16.650 965.075 16.930 965.445 ;
        RECT 16.720 959.470 16.860 965.075 ;
        RECT 16.660 959.150 16.920 959.470 ;
        RECT 608.680 959.150 608.940 959.470 ;
        RECT 608.740 749.770 608.880 959.150 ;
        RECT 609.390 749.770 609.670 750.000 ;
        RECT 608.740 749.630 609.670 749.770 ;
        RECT 609.390 746.000 609.670 749.630 ;
      LAYER via2 ;
        RECT 16.650 965.120 16.930 965.400 ;
      LAYER met3 ;
        RECT -4.800 965.410 2.400 965.860 ;
        RECT 16.625 965.410 16.955 965.425 ;
        RECT -4.800 965.110 16.955 965.410 ;
        RECT -4.800 964.660 2.400 965.110 ;
        RECT 16.625 965.095 16.955 965.110 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 459.610 747.900 459.930 747.960 ;
        RECT 459.610 747.760 483.070 747.900 ;
        RECT 459.610 747.700 459.930 747.760 ;
        RECT 429.800 747.420 432.700 747.560 ;
        RECT 17.090 746.880 17.410 746.940 ;
        RECT 429.800 746.880 429.940 747.420 ;
        RECT 17.090 746.740 429.940 746.880 ;
        RECT 432.560 746.880 432.700 747.420 ;
        RECT 459.610 747.020 459.930 747.280 ;
        RECT 459.700 746.880 459.840 747.020 ;
        RECT 432.560 746.740 459.840 746.880 ;
        RECT 482.930 746.880 483.070 747.760 ;
        RECT 612.790 747.220 613.110 747.280 ;
        RECT 572.860 747.080 613.110 747.220 ;
        RECT 572.860 746.880 573.000 747.080 ;
        RECT 612.790 747.020 613.110 747.080 ;
        RECT 482.930 746.740 573.000 746.880 ;
        RECT 17.090 746.680 17.410 746.740 ;
      LAYER via ;
        RECT 459.640 747.700 459.900 747.960 ;
        RECT 17.120 746.680 17.380 746.940 ;
        RECT 459.640 747.020 459.900 747.280 ;
        RECT 612.820 747.020 613.080 747.280 ;
      LAYER met2 ;
        RECT 459.640 747.670 459.900 747.990 ;
        RECT 459.700 747.310 459.840 747.670 ;
        RECT 459.640 746.990 459.900 747.310 ;
        RECT 612.820 747.050 613.080 747.310 ;
        RECT 613.530 747.050 613.810 750.000 ;
        RECT 612.820 746.990 613.810 747.050 ;
        RECT 17.120 746.650 17.380 746.970 ;
        RECT 612.880 746.910 613.810 746.990 ;
        RECT 17.180 714.525 17.320 746.650 ;
        RECT 613.530 746.000 613.810 746.910 ;
        RECT 17.110 714.155 17.390 714.525 ;
      LAYER via2 ;
        RECT 17.110 714.200 17.390 714.480 ;
      LAYER met3 ;
        RECT -4.800 714.490 2.400 714.940 ;
        RECT 17.085 714.490 17.415 714.505 ;
        RECT -4.800 714.190 17.415 714.490 ;
        RECT -4.800 713.740 2.400 714.190 ;
        RECT 17.085 714.175 17.415 714.190 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.390 753.680 19.710 753.740 ;
        RECT 616.930 753.680 617.250 753.740 ;
        RECT 19.390 753.540 617.250 753.680 ;
        RECT 19.390 753.480 19.710 753.540 ;
        RECT 616.930 753.480 617.250 753.540 ;
      LAYER via ;
        RECT 19.420 753.480 19.680 753.740 ;
        RECT 616.960 753.480 617.220 753.740 ;
      LAYER met2 ;
        RECT 19.420 753.450 19.680 753.770 ;
        RECT 616.960 753.450 617.220 753.770 ;
        RECT 19.480 463.605 19.620 753.450 ;
        RECT 617.020 749.770 617.160 753.450 ;
        RECT 617.670 749.770 617.950 750.000 ;
        RECT 617.020 749.630 617.950 749.770 ;
        RECT 617.670 746.000 617.950 749.630 ;
        RECT 19.410 463.235 19.690 463.605 ;
      LAYER via2 ;
        RECT 19.410 463.280 19.690 463.560 ;
      LAYER met3 ;
        RECT -4.800 463.570 2.400 464.020 ;
        RECT 19.385 463.570 19.715 463.585 ;
        RECT -4.800 463.270 19.715 463.570 ;
        RECT -4.800 462.820 2.400 463.270 ;
        RECT 19.385 463.255 19.715 463.270 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 753.000 18.330 753.060 ;
        RECT 621.070 753.000 621.390 753.060 ;
        RECT 18.010 752.860 621.390 753.000 ;
        RECT 18.010 752.800 18.330 752.860 ;
        RECT 621.070 752.800 621.390 752.860 ;
      LAYER via ;
        RECT 18.040 752.800 18.300 753.060 ;
        RECT 621.100 752.800 621.360 753.060 ;
      LAYER met2 ;
        RECT 18.040 752.770 18.300 753.090 ;
        RECT 621.100 752.770 621.360 753.090 ;
        RECT 18.100 212.685 18.240 752.770 ;
        RECT 621.160 749.770 621.300 752.770 ;
        RECT 621.810 749.770 622.090 750.000 ;
        RECT 621.160 749.630 622.090 749.770 ;
        RECT 621.810 746.000 622.090 749.630 ;
        RECT 18.030 212.315 18.310 212.685 ;
      LAYER via2 ;
        RECT 18.030 212.360 18.310 212.640 ;
      LAYER met3 ;
        RECT -4.800 212.650 2.400 213.100 ;
        RECT 18.005 212.650 18.335 212.665 ;
        RECT -4.800 212.350 18.335 212.650 ;
        RECT -4.800 211.900 2.400 212.350 ;
        RECT 18.005 212.335 18.335 212.350 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.590 752.320 442.910 752.380 ;
        RECT 2900.830 752.320 2901.150 752.380 ;
        RECT 442.590 752.180 2901.150 752.320 ;
        RECT 442.590 752.120 442.910 752.180 ;
        RECT 2900.830 752.120 2901.150 752.180 ;
      LAYER via ;
        RECT 442.620 752.120 442.880 752.380 ;
        RECT 2900.860 752.120 2901.120 752.380 ;
      LAYER met2 ;
        RECT 442.620 752.090 442.880 752.410 ;
        RECT 2900.860 752.090 2901.120 752.410 ;
        RECT 442.680 750.000 442.820 752.090 ;
        RECT 442.410 749.630 442.820 750.000 ;
        RECT 442.410 746.000 442.690 749.630 ;
        RECT 2900.920 743.085 2901.060 752.090 ;
        RECT 2900.850 742.715 2901.130 743.085 ;
      LAYER via2 ;
        RECT 2900.850 742.760 2901.130 743.040 ;
      LAYER met3 ;
        RECT 2900.825 743.050 2901.155 743.065 ;
        RECT 2917.600 743.050 2924.800 743.500 ;
        RECT 2900.825 742.750 2924.800 743.050 ;
        RECT 2900.825 742.735 2901.155 742.750 ;
        RECT 2917.600 742.300 2924.800 742.750 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 972.980 441.990 973.040 ;
        RECT 2900.830 972.980 2901.150 973.040 ;
        RECT 441.670 972.840 2901.150 972.980 ;
        RECT 441.670 972.780 441.990 972.840 ;
        RECT 2900.830 972.780 2901.150 972.840 ;
        RECT 441.670 801.280 441.990 801.340 ;
        RECT 447.190 801.280 447.510 801.340 ;
        RECT 441.670 801.140 447.510 801.280 ;
        RECT 441.670 801.080 441.990 801.140 ;
        RECT 447.190 801.080 447.510 801.140 ;
      LAYER via ;
        RECT 441.700 972.780 441.960 973.040 ;
        RECT 2900.860 972.780 2901.120 973.040 ;
        RECT 441.700 801.080 441.960 801.340 ;
        RECT 447.220 801.080 447.480 801.340 ;
      LAYER met2 ;
        RECT 2900.850 977.315 2901.130 977.685 ;
        RECT 2900.920 973.070 2901.060 977.315 ;
        RECT 441.700 972.750 441.960 973.070 ;
        RECT 2900.860 972.750 2901.120 973.070 ;
        RECT 441.760 801.370 441.900 972.750 ;
        RECT 441.700 801.050 441.960 801.370 ;
        RECT 447.220 801.050 447.480 801.370 ;
        RECT 447.280 749.770 447.420 801.050 ;
        RECT 447.930 749.770 448.210 750.000 ;
        RECT 447.280 749.630 448.210 749.770 ;
        RECT 447.930 746.000 448.210 749.630 ;
      LAYER via2 ;
        RECT 2900.850 977.360 2901.130 977.640 ;
      LAYER met3 ;
        RECT 2900.825 977.650 2901.155 977.665 ;
        RECT 2917.600 977.650 2924.800 978.100 ;
        RECT 2900.825 977.350 2924.800 977.650 ;
        RECT 2900.825 977.335 2901.155 977.350 ;
        RECT 2917.600 976.900 2924.800 977.350 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.950 1207.580 450.270 1207.640 ;
        RECT 2900.830 1207.580 2901.150 1207.640 ;
        RECT 449.950 1207.440 2901.150 1207.580 ;
        RECT 449.950 1207.380 450.270 1207.440 ;
        RECT 2900.830 1207.380 2901.150 1207.440 ;
        RECT 449.950 766.600 450.270 766.660 ;
        RECT 452.710 766.600 453.030 766.660 ;
        RECT 449.950 766.460 453.030 766.600 ;
        RECT 449.950 766.400 450.270 766.460 ;
        RECT 452.710 766.400 453.030 766.460 ;
      LAYER via ;
        RECT 449.980 1207.380 450.240 1207.640 ;
        RECT 2900.860 1207.380 2901.120 1207.640 ;
        RECT 449.980 766.400 450.240 766.660 ;
        RECT 452.740 766.400 453.000 766.660 ;
      LAYER met2 ;
        RECT 2900.850 1211.915 2901.130 1212.285 ;
        RECT 2900.920 1207.670 2901.060 1211.915 ;
        RECT 449.980 1207.350 450.240 1207.670 ;
        RECT 2900.860 1207.350 2901.120 1207.670 ;
        RECT 450.040 766.690 450.180 1207.350 ;
        RECT 449.980 766.370 450.240 766.690 ;
        RECT 452.740 766.370 453.000 766.690 ;
        RECT 452.800 749.770 452.940 766.370 ;
        RECT 453.450 749.770 453.730 750.000 ;
        RECT 452.800 749.630 453.730 749.770 ;
        RECT 453.450 746.000 453.730 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1211.960 2901.130 1212.240 ;
      LAYER met3 ;
        RECT 2900.825 1212.250 2901.155 1212.265 ;
        RECT 2917.600 1212.250 2924.800 1212.700 ;
        RECT 2900.825 1211.950 2924.800 1212.250 ;
        RECT 2900.825 1211.935 2901.155 1211.950 ;
        RECT 2917.600 1211.500 2924.800 1211.950 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.230 1442.180 458.550 1442.240 ;
        RECT 2900.830 1442.180 2901.150 1442.240 ;
        RECT 458.230 1442.040 2901.150 1442.180 ;
        RECT 458.230 1441.980 458.550 1442.040 ;
        RECT 2900.830 1441.980 2901.150 1442.040 ;
      LAYER via ;
        RECT 458.260 1441.980 458.520 1442.240 ;
        RECT 2900.860 1441.980 2901.120 1442.240 ;
      LAYER met2 ;
        RECT 2900.850 1446.515 2901.130 1446.885 ;
        RECT 2900.920 1442.270 2901.060 1446.515 ;
        RECT 458.260 1441.950 458.520 1442.270 ;
        RECT 2900.860 1441.950 2901.120 1442.270 ;
        RECT 458.320 749.770 458.460 1441.950 ;
        RECT 458.970 749.770 459.250 750.000 ;
        RECT 458.320 749.630 459.250 749.770 ;
        RECT 458.970 746.000 459.250 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1446.560 2901.130 1446.840 ;
      LAYER met3 ;
        RECT 2900.825 1446.850 2901.155 1446.865 ;
        RECT 2917.600 1446.850 2924.800 1447.300 ;
        RECT 2900.825 1446.550 2924.800 1446.850 ;
        RECT 2900.825 1446.535 2901.155 1446.550 ;
        RECT 2917.600 1446.100 2924.800 1446.550 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.210 1676.780 464.530 1676.840 ;
        RECT 2900.830 1676.780 2901.150 1676.840 ;
        RECT 464.210 1676.640 2901.150 1676.780 ;
        RECT 464.210 1676.580 464.530 1676.640 ;
        RECT 2900.830 1676.580 2901.150 1676.640 ;
      LAYER via ;
        RECT 464.240 1676.580 464.500 1676.840 ;
        RECT 2900.860 1676.580 2901.120 1676.840 ;
      LAYER met2 ;
        RECT 2900.850 1681.115 2901.130 1681.485 ;
        RECT 2900.920 1676.870 2901.060 1681.115 ;
        RECT 464.240 1676.550 464.500 1676.870 ;
        RECT 2900.860 1676.550 2901.120 1676.870 ;
        RECT 464.300 751.130 464.440 1676.550 ;
        RECT 464.300 750.990 464.670 751.130 ;
        RECT 464.530 750.000 464.670 750.990 ;
        RECT 464.490 746.000 464.770 750.000 ;
      LAYER via2 ;
        RECT 2900.850 1681.160 2901.130 1681.440 ;
      LAYER met3 ;
        RECT 2900.825 1681.450 2901.155 1681.465 ;
        RECT 2917.600 1681.450 2924.800 1681.900 ;
        RECT 2900.825 1681.150 2924.800 1681.450 ;
        RECT 2900.825 1681.135 2901.155 1681.150 ;
        RECT 2917.600 1680.700 2924.800 1681.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.730 1911.380 470.050 1911.440 ;
        RECT 2900.830 1911.380 2901.150 1911.440 ;
        RECT 469.730 1911.240 2901.150 1911.380 ;
        RECT 469.730 1911.180 470.050 1911.240 ;
        RECT 2900.830 1911.180 2901.150 1911.240 ;
      LAYER via ;
        RECT 469.760 1911.180 470.020 1911.440 ;
        RECT 2900.860 1911.180 2901.120 1911.440 ;
      LAYER met2 ;
        RECT 2900.850 1915.715 2901.130 1916.085 ;
        RECT 2900.920 1911.470 2901.060 1915.715 ;
        RECT 469.760 1911.150 470.020 1911.470 ;
        RECT 2900.860 1911.150 2901.120 1911.470 ;
        RECT 469.820 751.130 469.960 1911.150 ;
        RECT 469.820 750.990 470.190 751.130 ;
        RECT 470.050 750.000 470.190 750.990 ;
        RECT 470.010 746.000 470.290 750.000 ;
      LAYER via2 ;
        RECT 2900.850 1915.760 2901.130 1916.040 ;
      LAYER met3 ;
        RECT 2900.825 1916.050 2901.155 1916.065 ;
        RECT 2917.600 1916.050 2924.800 1916.500 ;
        RECT 2900.825 1915.750 2924.800 1916.050 ;
        RECT 2900.825 1915.735 2901.155 1915.750 ;
        RECT 2917.600 1915.300 2924.800 1915.750 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 473.410 2145.980 473.730 2146.040 ;
        RECT 2900.830 2145.980 2901.150 2146.040 ;
        RECT 473.410 2145.840 2901.150 2145.980 ;
        RECT 473.410 2145.780 473.730 2145.840 ;
        RECT 2900.830 2145.780 2901.150 2145.840 ;
      LAYER via ;
        RECT 473.440 2145.780 473.700 2146.040 ;
        RECT 2900.860 2145.780 2901.120 2146.040 ;
      LAYER met2 ;
        RECT 2900.850 2150.315 2901.130 2150.685 ;
        RECT 2900.920 2146.070 2901.060 2150.315 ;
        RECT 473.440 2145.750 473.700 2146.070 ;
        RECT 2900.860 2145.750 2901.120 2146.070 ;
        RECT 473.500 855.670 473.640 2145.750 ;
        RECT 473.500 855.530 475.020 855.670 ;
        RECT 474.880 749.770 475.020 855.530 ;
        RECT 475.530 749.770 475.810 750.000 ;
        RECT 474.880 749.630 475.810 749.770 ;
        RECT 475.530 746.000 475.810 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2150.360 2901.130 2150.640 ;
      LAYER met3 ;
        RECT 2900.825 2150.650 2901.155 2150.665 ;
        RECT 2917.600 2150.650 2924.800 2151.100 ;
        RECT 2900.825 2150.350 2924.800 2150.650 ;
        RECT 2900.825 2150.335 2901.155 2150.350 ;
        RECT 2917.600 2149.900 2924.800 2150.350 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 752.235 427.710 752.605 ;
        RECT 427.500 750.000 427.640 752.235 ;
        RECT 427.230 749.630 427.640 750.000 ;
        RECT 427.230 746.000 427.510 749.630 ;
      LAYER via2 ;
        RECT 427.430 752.280 427.710 752.560 ;
      LAYER met3 ;
        RECT 427.405 752.570 427.735 752.585 ;
        RECT 644.270 752.570 644.650 752.580 ;
        RECT 427.405 752.270 644.650 752.570 ;
        RECT 427.405 752.255 427.735 752.270 ;
        RECT 644.270 752.260 644.650 752.270 ;
        RECT 2917.600 195.650 2924.800 196.100 ;
        RECT 2916.710 195.350 2924.800 195.650 ;
        RECT 2916.710 194.970 2917.010 195.350 ;
        RECT 2917.600 194.970 2924.800 195.350 ;
        RECT 2916.710 194.900 2924.800 194.970 ;
        RECT 2916.710 194.670 2917.930 194.900 ;
        RECT 644.270 193.610 644.650 193.620 ;
        RECT 2917.630 193.610 2917.930 194.670 ;
        RECT 644.270 193.310 2917.930 193.610 ;
        RECT 644.270 193.300 644.650 193.310 ;
      LAYER via3 ;
        RECT 644.300 752.260 644.620 752.580 ;
        RECT 644.300 193.300 644.620 193.620 ;
      LAYER met4 ;
        RECT 644.295 752.255 644.625 752.585 ;
        RECT 644.310 193.625 644.610 752.255 ;
        RECT 644.295 193.295 644.625 193.625 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.930 2539.360 479.250 2539.420 ;
        RECT 2900.830 2539.360 2901.150 2539.420 ;
        RECT 478.930 2539.220 2901.150 2539.360 ;
        RECT 478.930 2539.160 479.250 2539.220 ;
        RECT 2900.830 2539.160 2901.150 2539.220 ;
      LAYER via ;
        RECT 478.960 2539.160 479.220 2539.420 ;
        RECT 2900.860 2539.160 2901.120 2539.420 ;
      LAYER met2 ;
        RECT 2900.850 2541.315 2901.130 2541.685 ;
        RECT 2900.920 2539.450 2901.060 2541.315 ;
        RECT 478.960 2539.130 479.220 2539.450 ;
        RECT 2900.860 2539.130 2901.120 2539.450 ;
        RECT 479.020 855.670 479.160 2539.130 ;
        RECT 479.020 855.530 481.920 855.670 ;
        RECT 481.780 749.770 481.920 855.530 ;
        RECT 482.430 749.770 482.710 750.000 ;
        RECT 481.780 749.630 482.710 749.770 ;
        RECT 482.430 746.000 482.710 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2541.360 2901.130 2541.640 ;
      LAYER met3 ;
        RECT 2900.825 2541.650 2901.155 2541.665 ;
        RECT 2917.600 2541.650 2924.800 2542.100 ;
        RECT 2900.825 2541.350 2924.800 2541.650 ;
        RECT 2900.825 2541.335 2901.155 2541.350 ;
        RECT 2917.600 2540.900 2924.800 2541.350 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.210 2773.960 487.530 2774.020 ;
        RECT 2900.830 2773.960 2901.150 2774.020 ;
        RECT 487.210 2773.820 2901.150 2773.960 ;
        RECT 487.210 2773.760 487.530 2773.820 ;
        RECT 2900.830 2773.760 2901.150 2773.820 ;
      LAYER via ;
        RECT 487.240 2773.760 487.500 2774.020 ;
        RECT 2900.860 2773.760 2901.120 2774.020 ;
      LAYER met2 ;
        RECT 2900.850 2775.915 2901.130 2776.285 ;
        RECT 2900.920 2774.050 2901.060 2775.915 ;
        RECT 487.240 2773.730 487.500 2774.050 ;
        RECT 2900.860 2773.730 2901.120 2774.050 ;
        RECT 487.300 749.770 487.440 2773.730 ;
        RECT 487.950 749.770 488.230 750.000 ;
        RECT 487.300 749.630 488.230 749.770 ;
        RECT 487.950 746.000 488.230 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2775.960 2901.130 2776.240 ;
      LAYER met3 ;
        RECT 2900.825 2776.250 2901.155 2776.265 ;
        RECT 2917.600 2776.250 2924.800 2776.700 ;
        RECT 2900.825 2775.950 2924.800 2776.250 ;
        RECT 2900.825 2775.935 2901.155 2775.950 ;
        RECT 2917.600 2775.500 2924.800 2775.950 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.730 3008.560 493.050 3008.620 ;
        RECT 2900.830 3008.560 2901.150 3008.620 ;
        RECT 492.730 3008.420 2901.150 3008.560 ;
        RECT 492.730 3008.360 493.050 3008.420 ;
        RECT 2900.830 3008.360 2901.150 3008.420 ;
      LAYER via ;
        RECT 492.760 3008.360 493.020 3008.620 ;
        RECT 2900.860 3008.360 2901.120 3008.620 ;
      LAYER met2 ;
        RECT 2900.850 3010.515 2901.130 3010.885 ;
        RECT 2900.920 3008.650 2901.060 3010.515 ;
        RECT 492.760 3008.330 493.020 3008.650 ;
        RECT 2900.860 3008.330 2901.120 3008.650 ;
        RECT 492.820 749.770 492.960 3008.330 ;
        RECT 493.470 749.770 493.750 750.000 ;
        RECT 492.820 749.630 493.750 749.770 ;
        RECT 493.470 746.000 493.750 749.630 ;
      LAYER via2 ;
        RECT 2900.850 3010.560 2901.130 3010.840 ;
      LAYER met3 ;
        RECT 2900.825 3010.850 2901.155 3010.865 ;
        RECT 2917.600 3010.850 2924.800 3011.300 ;
        RECT 2900.825 3010.550 2924.800 3010.850 ;
        RECT 2900.825 3010.535 2901.155 3010.550 ;
        RECT 2917.600 3010.100 2924.800 3010.550 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.250 3243.160 498.570 3243.220 ;
        RECT 2900.830 3243.160 2901.150 3243.220 ;
        RECT 498.250 3243.020 2901.150 3243.160 ;
        RECT 498.250 3242.960 498.570 3243.020 ;
        RECT 2900.830 3242.960 2901.150 3243.020 ;
      LAYER via ;
        RECT 498.280 3242.960 498.540 3243.220 ;
        RECT 2900.860 3242.960 2901.120 3243.220 ;
      LAYER met2 ;
        RECT 2900.850 3245.115 2901.130 3245.485 ;
        RECT 2900.920 3243.250 2901.060 3245.115 ;
        RECT 498.280 3242.930 498.540 3243.250 ;
        RECT 2900.860 3242.930 2901.120 3243.250 ;
        RECT 498.340 749.770 498.480 3242.930 ;
        RECT 498.990 749.770 499.270 750.000 ;
        RECT 498.340 749.630 499.270 749.770 ;
        RECT 498.990 746.000 499.270 749.630 ;
      LAYER via2 ;
        RECT 2900.850 3245.160 2901.130 3245.440 ;
      LAYER met3 ;
        RECT 2900.825 3245.450 2901.155 3245.465 ;
        RECT 2917.600 3245.450 2924.800 3245.900 ;
        RECT 2900.825 3245.150 2924.800 3245.450 ;
        RECT 2900.825 3245.135 2901.155 3245.150 ;
        RECT 2917.600 3244.700 2924.800 3245.150 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 3477.760 504.550 3477.820 ;
        RECT 2900.830 3477.760 2901.150 3477.820 ;
        RECT 504.230 3477.620 2901.150 3477.760 ;
        RECT 504.230 3477.560 504.550 3477.620 ;
        RECT 2900.830 3477.560 2901.150 3477.620 ;
      LAYER via ;
        RECT 504.260 3477.560 504.520 3477.820 ;
        RECT 2900.860 3477.560 2901.120 3477.820 ;
      LAYER met2 ;
        RECT 2900.850 3479.715 2901.130 3480.085 ;
        RECT 2900.920 3477.850 2901.060 3479.715 ;
        RECT 504.260 3477.530 504.520 3477.850 ;
        RECT 2900.860 3477.530 2901.120 3477.850 ;
        RECT 504.320 751.130 504.460 3477.530 ;
        RECT 504.320 750.990 504.690 751.130 ;
        RECT 504.550 750.000 504.690 750.990 ;
        RECT 504.510 746.000 504.790 750.000 ;
      LAYER via2 ;
        RECT 2900.850 3479.760 2901.130 3480.040 ;
      LAYER met3 ;
        RECT 2900.825 3480.050 2901.155 3480.065 ;
        RECT 2917.600 3480.050 2924.800 3480.500 ;
        RECT 2900.825 3479.750 2924.800 3480.050 ;
        RECT 2900.825 3479.735 2901.155 3479.750 ;
        RECT 2917.600 3479.300 2924.800 3479.750 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.290 776.120 509.610 776.180 ;
        RECT 2642.770 776.120 2643.090 776.180 ;
        RECT 509.290 775.980 2643.090 776.120 ;
        RECT 509.290 775.920 509.610 775.980 ;
        RECT 2642.770 775.920 2643.090 775.980 ;
      LAYER via ;
        RECT 509.320 775.920 509.580 776.180 ;
        RECT 2642.800 775.920 2643.060 776.180 ;
      LAYER met2 ;
        RECT 2642.860 3517.910 2648.060 3518.050 ;
        RECT 2642.860 776.210 2643.000 3517.910 ;
        RECT 2647.920 3517.370 2648.060 3517.910 ;
        RECT 2648.630 3517.600 2649.190 3524.800 ;
        RECT 2648.840 3517.370 2648.980 3517.600 ;
        RECT 2647.920 3517.230 2648.980 3517.370 ;
        RECT 509.320 775.890 509.580 776.210 ;
        RECT 2642.800 775.890 2643.060 776.210 ;
        RECT 509.380 749.770 509.520 775.890 ;
        RECT 510.030 749.770 510.310 750.000 ;
        RECT 509.380 749.630 510.310 749.770 ;
        RECT 510.030 746.000 510.310 749.630 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2318.470 3515.160 2318.790 3515.220 ;
        RECT 2324.450 3515.160 2324.770 3515.220 ;
        RECT 2318.470 3515.020 2324.770 3515.160 ;
        RECT 2318.470 3514.960 2318.790 3515.020 ;
        RECT 2324.450 3514.960 2324.770 3515.020 ;
        RECT 514.810 776.460 515.130 776.520 ;
        RECT 2318.470 776.460 2318.790 776.520 ;
        RECT 514.810 776.320 2318.790 776.460 ;
        RECT 514.810 776.260 515.130 776.320 ;
        RECT 2318.470 776.260 2318.790 776.320 ;
      LAYER via ;
        RECT 2318.500 3514.960 2318.760 3515.220 ;
        RECT 2324.480 3514.960 2324.740 3515.220 ;
        RECT 514.840 776.260 515.100 776.520 ;
        RECT 2318.500 776.260 2318.760 776.520 ;
      LAYER met2 ;
        RECT 2324.330 3517.600 2324.890 3524.800 ;
        RECT 2324.540 3515.250 2324.680 3517.600 ;
        RECT 2318.500 3514.930 2318.760 3515.250 ;
        RECT 2324.480 3514.930 2324.740 3515.250 ;
        RECT 2318.560 776.550 2318.700 3514.930 ;
        RECT 514.840 776.230 515.100 776.550 ;
        RECT 2318.500 776.230 2318.760 776.550 ;
        RECT 514.900 749.770 515.040 776.230 ;
        RECT 515.550 749.770 515.830 750.000 ;
        RECT 514.900 749.630 515.830 749.770 ;
        RECT 515.550 746.000 515.830 749.630 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.330 776.800 520.650 776.860 ;
        RECT 1994.170 776.800 1994.490 776.860 ;
        RECT 520.330 776.660 1994.490 776.800 ;
        RECT 520.330 776.600 520.650 776.660 ;
        RECT 1994.170 776.600 1994.490 776.660 ;
      LAYER via ;
        RECT 520.360 776.600 520.620 776.860 ;
        RECT 1994.200 776.600 1994.460 776.860 ;
      LAYER met2 ;
        RECT 1994.260 3517.910 1999.460 3518.050 ;
        RECT 1994.260 776.890 1994.400 3517.910 ;
        RECT 1999.320 3517.370 1999.460 3517.910 ;
        RECT 2000.030 3517.600 2000.590 3524.800 ;
        RECT 2000.240 3517.370 2000.380 3517.600 ;
        RECT 1999.320 3517.230 2000.380 3517.370 ;
        RECT 520.360 776.570 520.620 776.890 ;
        RECT 1994.200 776.570 1994.460 776.890 ;
        RECT 520.420 749.770 520.560 776.570 ;
        RECT 521.070 749.770 521.350 750.000 ;
        RECT 520.420 749.630 521.350 749.770 ;
        RECT 521.070 746.000 521.350 749.630 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1669.870 3515.160 1670.190 3515.220 ;
        RECT 1675.850 3515.160 1676.170 3515.220 ;
        RECT 1669.870 3515.020 1676.170 3515.160 ;
        RECT 1669.870 3514.960 1670.190 3515.020 ;
        RECT 1675.850 3514.960 1676.170 3515.020 ;
        RECT 525.390 783.600 525.710 783.660 ;
        RECT 1669.870 783.600 1670.190 783.660 ;
        RECT 525.390 783.460 1670.190 783.600 ;
        RECT 525.390 783.400 525.710 783.460 ;
        RECT 1669.870 783.400 1670.190 783.460 ;
      LAYER via ;
        RECT 1669.900 3514.960 1670.160 3515.220 ;
        RECT 1675.880 3514.960 1676.140 3515.220 ;
        RECT 525.420 783.400 525.680 783.660 ;
        RECT 1669.900 783.400 1670.160 783.660 ;
      LAYER met2 ;
        RECT 1675.730 3517.600 1676.290 3524.800 ;
        RECT 1675.940 3515.250 1676.080 3517.600 ;
        RECT 1669.900 3514.930 1670.160 3515.250 ;
        RECT 1675.880 3514.930 1676.140 3515.250 ;
        RECT 1669.960 783.690 1670.100 3514.930 ;
        RECT 525.420 783.370 525.680 783.690 ;
        RECT 1669.900 783.370 1670.160 783.690 ;
        RECT 525.480 759.070 525.620 783.370 ;
        RECT 525.480 758.930 526.080 759.070 ;
        RECT 525.940 749.770 526.080 758.930 ;
        RECT 526.590 749.770 526.870 750.000 ;
        RECT 525.940 749.630 526.870 749.770 ;
        RECT 526.590 746.000 526.870 749.630 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 783.940 532.150 784.000 ;
        RECT 1345.570 783.940 1345.890 784.000 ;
        RECT 531.830 783.800 1345.890 783.940 ;
        RECT 531.830 783.740 532.150 783.800 ;
        RECT 1345.570 783.740 1345.890 783.800 ;
      LAYER via ;
        RECT 531.860 783.740 532.120 784.000 ;
        RECT 1345.600 783.740 1345.860 784.000 ;
      LAYER met2 ;
        RECT 1345.660 3517.910 1350.860 3518.050 ;
        RECT 1345.660 784.030 1345.800 3517.910 ;
        RECT 1350.720 3517.370 1350.860 3517.910 ;
        RECT 1351.430 3517.600 1351.990 3524.800 ;
        RECT 1351.640 3517.370 1351.780 3517.600 ;
        RECT 1350.720 3517.230 1351.780 3517.370 ;
        RECT 531.860 783.710 532.120 784.030 ;
        RECT 1345.600 783.710 1345.860 784.030 ;
        RECT 531.920 751.130 532.060 783.710 ;
        RECT 531.920 750.990 532.290 751.130 ;
        RECT 532.150 750.000 532.290 750.990 ;
        RECT 532.110 746.000 532.390 750.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 433.390 747.560 433.710 747.620 ;
        RECT 433.390 747.420 460.300 747.560 ;
        RECT 433.390 747.360 433.710 747.420 ;
        RECT 460.160 746.200 460.300 747.420 ;
        RECT 2902.670 746.200 2902.990 746.260 ;
        RECT 460.160 746.060 2902.990 746.200 ;
        RECT 2902.670 746.000 2902.990 746.060 ;
      LAYER via ;
        RECT 433.420 747.360 433.680 747.620 ;
        RECT 2902.700 746.000 2902.960 746.260 ;
      LAYER met2 ;
        RECT 432.750 747.730 433.030 750.000 ;
        RECT 432.750 747.650 433.620 747.730 ;
        RECT 432.750 747.590 433.680 747.650 ;
        RECT 432.750 746.000 433.030 747.590 ;
        RECT 433.420 747.330 433.680 747.590 ;
        RECT 2902.700 745.970 2902.960 746.290 ;
        RECT 2902.760 430.285 2902.900 745.970 ;
        RECT 2902.690 429.915 2902.970 430.285 ;
      LAYER via2 ;
        RECT 2902.690 429.960 2902.970 430.240 ;
      LAYER met3 ;
        RECT 2902.665 430.250 2902.995 430.265 ;
        RECT 2917.600 430.250 2924.800 430.700 ;
        RECT 2902.665 429.950 2924.800 430.250 ;
        RECT 2902.665 429.935 2902.995 429.950 ;
        RECT 2917.600 429.500 2924.800 429.950 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.270 3515.160 1021.590 3515.220 ;
        RECT 1027.250 3515.160 1027.570 3515.220 ;
        RECT 1021.270 3515.020 1027.570 3515.160 ;
        RECT 1021.270 3514.960 1021.590 3515.020 ;
        RECT 1027.250 3514.960 1027.570 3515.020 ;
        RECT 536.890 784.620 537.210 784.680 ;
        RECT 1021.270 784.620 1021.590 784.680 ;
        RECT 536.890 784.480 1021.590 784.620 ;
        RECT 536.890 784.420 537.210 784.480 ;
        RECT 1021.270 784.420 1021.590 784.480 ;
      LAYER via ;
        RECT 1021.300 3514.960 1021.560 3515.220 ;
        RECT 1027.280 3514.960 1027.540 3515.220 ;
        RECT 536.920 784.420 537.180 784.680 ;
        RECT 1021.300 784.420 1021.560 784.680 ;
      LAYER met2 ;
        RECT 1027.130 3517.600 1027.690 3524.800 ;
        RECT 1027.340 3515.250 1027.480 3517.600 ;
        RECT 1021.300 3514.930 1021.560 3515.250 ;
        RECT 1027.280 3514.930 1027.540 3515.250 ;
        RECT 1021.360 784.710 1021.500 3514.930 ;
        RECT 536.920 784.390 537.180 784.710 ;
        RECT 1021.300 784.390 1021.560 784.710 ;
        RECT 536.980 749.770 537.120 784.390 ;
        RECT 537.630 749.770 537.910 750.000 ;
        RECT 536.980 749.630 537.910 749.770 ;
        RECT 537.630 746.000 537.910 749.630 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 542.410 785.300 542.730 785.360 ;
        RECT 696.970 785.300 697.290 785.360 ;
        RECT 542.410 785.160 697.290 785.300 ;
        RECT 542.410 785.100 542.730 785.160 ;
        RECT 696.970 785.100 697.290 785.160 ;
      LAYER via ;
        RECT 542.440 785.100 542.700 785.360 ;
        RECT 697.000 785.100 697.260 785.360 ;
      LAYER met2 ;
        RECT 697.060 3517.910 702.260 3518.050 ;
        RECT 697.060 785.390 697.200 3517.910 ;
        RECT 702.120 3517.370 702.260 3517.910 ;
        RECT 702.830 3517.600 703.390 3524.800 ;
        RECT 703.040 3517.370 703.180 3517.600 ;
        RECT 702.120 3517.230 703.180 3517.370 ;
        RECT 542.440 785.070 542.700 785.390 ;
        RECT 697.000 785.070 697.260 785.390 ;
        RECT 542.500 749.770 542.640 785.070 ;
        RECT 543.150 749.770 543.430 750.000 ;
        RECT 542.500 749.630 543.430 749.770 ;
        RECT 543.150 746.000 543.430 749.630 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 3515.160 372.990 3515.220 ;
        RECT 378.650 3515.160 378.970 3515.220 ;
        RECT 372.670 3515.020 378.970 3515.160 ;
        RECT 372.670 3514.960 372.990 3515.020 ;
        RECT 378.650 3514.960 378.970 3515.020 ;
        RECT 372.670 784.960 372.990 785.020 ;
        RECT 548.390 784.960 548.710 785.020 ;
        RECT 372.670 784.820 548.710 784.960 ;
        RECT 372.670 784.760 372.990 784.820 ;
        RECT 548.390 784.760 548.710 784.820 ;
      LAYER via ;
        RECT 372.700 3514.960 372.960 3515.220 ;
        RECT 378.680 3514.960 378.940 3515.220 ;
        RECT 372.700 784.760 372.960 785.020 ;
        RECT 548.420 784.760 548.680 785.020 ;
      LAYER met2 ;
        RECT 378.530 3517.600 379.090 3524.800 ;
        RECT 378.740 3515.250 378.880 3517.600 ;
        RECT 372.700 3514.930 372.960 3515.250 ;
        RECT 378.680 3514.930 378.940 3515.250 ;
        RECT 372.760 785.050 372.900 3514.930 ;
        RECT 372.700 784.730 372.960 785.050 ;
        RECT 548.420 784.730 548.680 785.050 ;
        RECT 548.480 751.130 548.620 784.730 ;
        RECT 548.480 750.990 548.850 751.130 ;
        RECT 548.710 750.000 548.850 750.990 ;
        RECT 548.670 746.000 548.950 750.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 48.370 784.280 48.690 784.340 ;
        RECT 553.450 784.280 553.770 784.340 ;
        RECT 48.370 784.140 553.770 784.280 ;
        RECT 48.370 784.080 48.690 784.140 ;
        RECT 553.450 784.080 553.770 784.140 ;
      LAYER via ;
        RECT 48.400 784.080 48.660 784.340 ;
        RECT 553.480 784.080 553.740 784.340 ;
      LAYER met2 ;
        RECT 48.460 3517.910 53.660 3518.050 ;
        RECT 48.460 784.370 48.600 3517.910 ;
        RECT 53.520 3517.370 53.660 3517.910 ;
        RECT 54.230 3517.600 54.790 3524.800 ;
        RECT 54.440 3517.370 54.580 3517.600 ;
        RECT 53.520 3517.230 54.580 3517.370 ;
        RECT 48.400 784.050 48.660 784.370 ;
        RECT 553.480 784.050 553.740 784.370 ;
        RECT 553.540 749.770 553.680 784.050 ;
        RECT 554.190 749.770 554.470 750.000 ;
        RECT 553.540 749.630 554.470 749.770 ;
        RECT 554.190 746.000 554.470 749.630 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3305.380 17.410 3305.440 ;
        RECT 559.430 3305.380 559.750 3305.440 ;
        RECT 17.090 3305.240 559.750 3305.380 ;
        RECT 17.090 3305.180 17.410 3305.240 ;
        RECT 559.430 3305.180 559.750 3305.240 ;
      LAYER via ;
        RECT 17.120 3305.180 17.380 3305.440 ;
        RECT 559.460 3305.180 559.720 3305.440 ;
      LAYER met2 ;
        RECT 17.110 3306.995 17.390 3307.365 ;
        RECT 17.180 3305.470 17.320 3306.995 ;
        RECT 17.120 3305.150 17.380 3305.470 ;
        RECT 559.460 3305.150 559.720 3305.470 ;
        RECT 559.520 751.130 559.660 3305.150 ;
        RECT 559.520 750.990 559.890 751.130 ;
        RECT 559.750 750.000 559.890 750.990 ;
        RECT 559.710 746.000 559.990 750.000 ;
      LAYER via2 ;
        RECT 17.110 3307.040 17.390 3307.320 ;
      LAYER met3 ;
        RECT -4.800 3307.330 2.400 3307.780 ;
        RECT 17.085 3307.330 17.415 3307.345 ;
        RECT -4.800 3307.030 17.415 3307.330 ;
        RECT -4.800 3306.580 2.400 3307.030 ;
        RECT 17.085 3307.015 17.415 3307.030 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 555.290 3050.040 555.610 3050.100 ;
        RECT 17.090 3049.900 555.610 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 555.290 3049.840 555.610 3049.900 ;
        RECT 555.290 765.920 555.610 765.980 ;
        RECT 564.490 765.920 564.810 765.980 ;
        RECT 555.290 765.780 564.810 765.920 ;
        RECT 555.290 765.720 555.610 765.780 ;
        RECT 564.490 765.720 564.810 765.780 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 555.320 3049.840 555.580 3050.100 ;
        RECT 555.320 765.720 555.580 765.980 ;
        RECT 564.520 765.720 564.780 765.980 ;
      LAYER met2 ;
        RECT 17.110 3056.075 17.390 3056.445 ;
        RECT 17.180 3050.130 17.320 3056.075 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 555.320 3049.810 555.580 3050.130 ;
        RECT 555.380 766.010 555.520 3049.810 ;
        RECT 555.320 765.690 555.580 766.010 ;
        RECT 564.520 765.690 564.780 766.010 ;
        RECT 564.580 749.770 564.720 765.690 ;
        RECT 565.230 749.770 565.510 750.000 ;
        RECT 564.580 749.630 565.510 749.770 ;
        RECT 565.230 746.000 565.510 749.630 ;
      LAYER via2 ;
        RECT 17.110 3056.120 17.390 3056.400 ;
      LAYER met3 ;
        RECT -4.800 3056.410 2.400 3056.860 ;
        RECT 17.085 3056.410 17.415 3056.425 ;
        RECT -4.800 3056.110 17.415 3056.410 ;
        RECT -4.800 3055.660 2.400 3056.110 ;
        RECT 17.085 3056.095 17.415 3056.110 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2801.500 15.570 2801.560 ;
        RECT 562.190 2801.500 562.510 2801.560 ;
        RECT 15.250 2801.360 562.510 2801.500 ;
        RECT 15.250 2801.300 15.570 2801.360 ;
        RECT 562.190 2801.300 562.510 2801.360 ;
        RECT 562.190 759.460 562.510 759.520 ;
        RECT 570.010 759.460 570.330 759.520 ;
        RECT 562.190 759.320 570.330 759.460 ;
        RECT 562.190 759.260 562.510 759.320 ;
        RECT 570.010 759.260 570.330 759.320 ;
      LAYER via ;
        RECT 15.280 2801.300 15.540 2801.560 ;
        RECT 562.220 2801.300 562.480 2801.560 ;
        RECT 562.220 759.260 562.480 759.520 ;
        RECT 570.040 759.260 570.300 759.520 ;
      LAYER met2 ;
        RECT 15.270 2805.155 15.550 2805.525 ;
        RECT 15.340 2801.590 15.480 2805.155 ;
        RECT 15.280 2801.270 15.540 2801.590 ;
        RECT 562.220 2801.270 562.480 2801.590 ;
        RECT 562.280 759.550 562.420 2801.270 ;
        RECT 562.220 759.230 562.480 759.550 ;
        RECT 570.040 759.230 570.300 759.550 ;
        RECT 570.100 749.770 570.240 759.230 ;
        RECT 570.750 749.770 571.030 750.000 ;
        RECT 570.100 749.630 571.030 749.770 ;
        RECT 570.750 746.000 571.030 749.630 ;
      LAYER via2 ;
        RECT 15.270 2805.200 15.550 2805.480 ;
      LAYER met3 ;
        RECT -4.800 2805.490 2.400 2805.940 ;
        RECT 15.245 2805.490 15.575 2805.505 ;
        RECT -4.800 2805.190 15.575 2805.490 ;
        RECT -4.800 2804.740 2.400 2805.190 ;
        RECT 15.245 2805.175 15.575 2805.190 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2553.300 16.950 2553.360 ;
        RECT 562.650 2553.300 562.970 2553.360 ;
        RECT 16.630 2553.160 562.970 2553.300 ;
        RECT 16.630 2553.100 16.950 2553.160 ;
        RECT 562.650 2553.100 562.970 2553.160 ;
        RECT 562.650 759.120 562.970 759.180 ;
        RECT 575.070 759.120 575.390 759.180 ;
        RECT 562.650 758.980 575.390 759.120 ;
        RECT 562.650 758.920 562.970 758.980 ;
        RECT 575.070 758.920 575.390 758.980 ;
      LAYER via ;
        RECT 16.660 2553.100 16.920 2553.360 ;
        RECT 562.680 2553.100 562.940 2553.360 ;
        RECT 562.680 758.920 562.940 759.180 ;
        RECT 575.100 758.920 575.360 759.180 ;
      LAYER met2 ;
        RECT 16.650 2554.235 16.930 2554.605 ;
        RECT 16.720 2553.390 16.860 2554.235 ;
        RECT 16.660 2553.070 16.920 2553.390 ;
        RECT 562.680 2553.070 562.940 2553.390 ;
        RECT 562.740 759.210 562.880 2553.070 ;
        RECT 562.680 758.890 562.940 759.210 ;
        RECT 575.100 758.890 575.360 759.210 ;
        RECT 575.160 752.490 575.300 758.890 ;
        RECT 575.160 752.350 575.760 752.490 ;
        RECT 575.620 749.770 575.760 752.350 ;
        RECT 576.270 749.770 576.550 750.000 ;
        RECT 575.620 749.630 576.550 749.770 ;
        RECT 576.270 746.000 576.550 749.630 ;
      LAYER via2 ;
        RECT 16.650 2554.280 16.930 2554.560 ;
      LAYER met3 ;
        RECT -4.800 2554.570 2.400 2555.020 ;
        RECT 16.625 2554.570 16.955 2554.585 ;
        RECT -4.800 2554.270 16.955 2554.570 ;
        RECT -4.800 2553.820 2.400 2554.270 ;
        RECT 16.625 2554.255 16.955 2554.270 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2297.960 16.030 2298.020 ;
        RECT 569.090 2297.960 569.410 2298.020 ;
        RECT 15.710 2297.820 569.410 2297.960 ;
        RECT 15.710 2297.760 16.030 2297.820 ;
        RECT 569.090 2297.760 569.410 2297.820 ;
        RECT 569.090 765.920 569.410 765.980 ;
        RECT 581.510 765.920 581.830 765.980 ;
        RECT 569.090 765.780 581.830 765.920 ;
        RECT 569.090 765.720 569.410 765.780 ;
        RECT 581.510 765.720 581.830 765.780 ;
      LAYER via ;
        RECT 15.740 2297.760 16.000 2298.020 ;
        RECT 569.120 2297.760 569.380 2298.020 ;
        RECT 569.120 765.720 569.380 765.980 ;
        RECT 581.540 765.720 581.800 765.980 ;
      LAYER met2 ;
        RECT 15.730 2303.315 16.010 2303.685 ;
        RECT 15.800 2298.050 15.940 2303.315 ;
        RECT 15.740 2297.730 16.000 2298.050 ;
        RECT 569.120 2297.730 569.380 2298.050 ;
        RECT 569.180 766.010 569.320 2297.730 ;
        RECT 569.120 765.690 569.380 766.010 ;
        RECT 581.540 765.690 581.800 766.010 ;
        RECT 581.600 751.130 581.740 765.690 ;
        RECT 581.600 750.990 581.970 751.130 ;
        RECT 581.830 750.000 581.970 750.990 ;
        RECT 581.790 746.000 582.070 750.000 ;
      LAYER via2 ;
        RECT 15.730 2303.360 16.010 2303.640 ;
      LAYER met3 ;
        RECT -4.800 2303.650 2.400 2304.100 ;
        RECT 15.705 2303.650 16.035 2303.665 ;
        RECT -4.800 2303.350 16.035 2303.650 ;
        RECT -4.800 2302.900 2.400 2303.350 ;
        RECT 15.705 2303.335 16.035 2303.350 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2049.420 16.950 2049.480 ;
        RECT 569.550 2049.420 569.870 2049.480 ;
        RECT 16.630 2049.280 569.870 2049.420 ;
        RECT 16.630 2049.220 16.950 2049.280 ;
        RECT 569.550 2049.220 569.870 2049.280 ;
        RECT 569.550 779.520 569.870 779.580 ;
        RECT 587.490 779.520 587.810 779.580 ;
        RECT 569.550 779.380 587.810 779.520 ;
        RECT 569.550 779.320 569.870 779.380 ;
        RECT 587.490 779.320 587.810 779.380 ;
      LAYER via ;
        RECT 16.660 2049.220 16.920 2049.480 ;
        RECT 569.580 2049.220 569.840 2049.480 ;
        RECT 569.580 779.320 569.840 779.580 ;
        RECT 587.520 779.320 587.780 779.580 ;
      LAYER met2 ;
        RECT 16.650 2052.395 16.930 2052.765 ;
        RECT 16.720 2049.510 16.860 2052.395 ;
        RECT 16.660 2049.190 16.920 2049.510 ;
        RECT 569.580 2049.190 569.840 2049.510 ;
        RECT 569.640 779.610 569.780 2049.190 ;
        RECT 569.580 779.290 569.840 779.610 ;
        RECT 587.520 779.290 587.780 779.610 ;
        RECT 587.580 750.000 587.720 779.290 ;
        RECT 587.310 749.630 587.720 750.000 ;
        RECT 587.310 746.000 587.590 749.630 ;
      LAYER via2 ;
        RECT 16.650 2052.440 16.930 2052.720 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 16.625 2052.730 16.955 2052.745 ;
        RECT -4.800 2052.430 16.955 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 16.625 2052.415 16.955 2052.430 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.910 754.020 439.230 754.080 ;
        RECT 644.990 754.020 645.310 754.080 ;
        RECT 438.910 753.880 645.310 754.020 ;
        RECT 438.910 753.820 439.230 753.880 ;
        RECT 644.990 753.820 645.310 753.880 ;
        RECT 644.990 669.360 645.310 669.420 ;
        RECT 2899.910 669.360 2900.230 669.420 ;
        RECT 644.990 669.220 2900.230 669.360 ;
        RECT 644.990 669.160 645.310 669.220 ;
        RECT 2899.910 669.160 2900.230 669.220 ;
      LAYER via ;
        RECT 438.940 753.820 439.200 754.080 ;
        RECT 645.020 753.820 645.280 754.080 ;
        RECT 645.020 669.160 645.280 669.420 ;
        RECT 2899.940 669.160 2900.200 669.420 ;
      LAYER met2 ;
        RECT 438.940 753.790 439.200 754.110 ;
        RECT 645.020 753.790 645.280 754.110 ;
        RECT 438.270 749.770 438.550 750.000 ;
        RECT 439.000 749.770 439.140 753.790 ;
        RECT 438.270 749.630 439.140 749.770 ;
        RECT 438.270 746.000 438.550 749.630 ;
        RECT 645.080 669.450 645.220 753.790 ;
        RECT 645.020 669.130 645.280 669.450 ;
        RECT 2899.940 669.130 2900.200 669.450 ;
        RECT 2900.000 664.885 2900.140 669.130 ;
        RECT 2899.930 664.515 2900.210 664.885 ;
      LAYER via2 ;
        RECT 2899.930 664.560 2900.210 664.840 ;
      LAYER met3 ;
        RECT 2899.905 664.850 2900.235 664.865 ;
        RECT 2917.600 664.850 2924.800 665.300 ;
        RECT 2899.905 664.550 2924.800 664.850 ;
        RECT 2899.905 664.535 2900.235 664.550 ;
        RECT 2917.600 664.100 2924.800 664.550 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1801.220 16.950 1801.280 ;
        RECT 575.990 1801.220 576.310 1801.280 ;
        RECT 16.630 1801.080 576.310 1801.220 ;
        RECT 16.630 1801.020 16.950 1801.080 ;
        RECT 575.990 1801.020 576.310 1801.080 ;
        RECT 575.990 765.580 576.310 765.640 ;
        RECT 592.090 765.580 592.410 765.640 ;
        RECT 575.990 765.440 592.410 765.580 ;
        RECT 575.990 765.380 576.310 765.440 ;
        RECT 592.090 765.380 592.410 765.440 ;
      LAYER via ;
        RECT 16.660 1801.020 16.920 1801.280 ;
        RECT 576.020 1801.020 576.280 1801.280 ;
        RECT 576.020 765.380 576.280 765.640 ;
        RECT 592.120 765.380 592.380 765.640 ;
      LAYER met2 ;
        RECT 16.650 1801.475 16.930 1801.845 ;
        RECT 16.720 1801.310 16.860 1801.475 ;
        RECT 16.660 1800.990 16.920 1801.310 ;
        RECT 576.020 1800.990 576.280 1801.310 ;
        RECT 576.080 765.670 576.220 1800.990 ;
        RECT 576.020 765.350 576.280 765.670 ;
        RECT 592.120 765.350 592.380 765.670 ;
        RECT 592.180 749.770 592.320 765.350 ;
        RECT 592.830 749.770 593.110 750.000 ;
        RECT 592.180 749.630 593.110 749.770 ;
        RECT 592.830 746.000 593.110 749.630 ;
      LAYER via2 ;
        RECT 16.650 1801.520 16.930 1801.800 ;
      LAYER met3 ;
        RECT -4.800 1801.810 2.400 1802.260 ;
        RECT 16.625 1801.810 16.955 1801.825 ;
        RECT -4.800 1801.510 16.955 1801.810 ;
        RECT -4.800 1801.060 2.400 1801.510 ;
        RECT 16.625 1801.495 16.955 1801.510 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.880 16.950 1545.940 ;
        RECT 598.070 1545.880 598.390 1545.940 ;
        RECT 16.630 1545.740 598.390 1545.880 ;
        RECT 16.630 1545.680 16.950 1545.740 ;
        RECT 598.070 1545.680 598.390 1545.740 ;
      LAYER via ;
        RECT 16.660 1545.680 16.920 1545.940 ;
        RECT 598.100 1545.680 598.360 1545.940 ;
      LAYER met2 ;
        RECT 16.650 1550.555 16.930 1550.925 ;
        RECT 16.720 1545.970 16.860 1550.555 ;
        RECT 16.660 1545.650 16.920 1545.970 ;
        RECT 598.100 1545.650 598.360 1545.970 ;
        RECT 598.160 751.130 598.300 1545.650 ;
        RECT 598.160 750.990 598.530 751.130 ;
        RECT 598.390 750.000 598.530 750.990 ;
        RECT 598.350 746.000 598.630 750.000 ;
      LAYER via2 ;
        RECT 16.650 1550.600 16.930 1550.880 ;
      LAYER met3 ;
        RECT -4.800 1550.890 2.400 1551.340 ;
        RECT 16.625 1550.890 16.955 1550.905 ;
        RECT -4.800 1550.590 16.955 1550.890 ;
        RECT -4.800 1550.140 2.400 1550.590 ;
        RECT 16.625 1550.575 16.955 1550.590 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.790 1297.340 15.110 1297.400 ;
        RECT 602.210 1297.340 602.530 1297.400 ;
        RECT 14.790 1297.200 602.530 1297.340 ;
        RECT 14.790 1297.140 15.110 1297.200 ;
        RECT 602.210 1297.140 602.530 1297.200 ;
      LAYER via ;
        RECT 14.820 1297.140 15.080 1297.400 ;
        RECT 602.240 1297.140 602.500 1297.400 ;
      LAYER met2 ;
        RECT 14.810 1299.635 15.090 1300.005 ;
        RECT 14.880 1297.430 15.020 1299.635 ;
        RECT 14.820 1297.110 15.080 1297.430 ;
        RECT 602.240 1297.110 602.500 1297.430 ;
        RECT 602.300 751.130 602.440 1297.110 ;
        RECT 602.300 750.990 602.670 751.130 ;
        RECT 602.530 750.000 602.670 750.990 ;
        RECT 602.490 746.000 602.770 750.000 ;
      LAYER via2 ;
        RECT 14.810 1299.680 15.090 1299.960 ;
      LAYER met3 ;
        RECT -4.800 1299.970 2.400 1300.420 ;
        RECT 14.785 1299.970 15.115 1299.985 ;
        RECT -4.800 1299.670 15.115 1299.970 ;
        RECT -4.800 1299.220 2.400 1299.670 ;
        RECT 14.785 1299.655 15.115 1299.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1049.140 16.950 1049.200 ;
        RECT 582.890 1049.140 583.210 1049.200 ;
        RECT 16.630 1049.000 583.210 1049.140 ;
        RECT 16.630 1048.940 16.950 1049.000 ;
        RECT 582.890 1048.940 583.210 1049.000 ;
        RECT 582.890 765.240 583.210 765.300 ;
        RECT 605.890 765.240 606.210 765.300 ;
        RECT 582.890 765.100 606.210 765.240 ;
        RECT 582.890 765.040 583.210 765.100 ;
        RECT 605.890 765.040 606.210 765.100 ;
      LAYER via ;
        RECT 16.660 1048.940 16.920 1049.200 ;
        RECT 582.920 1048.940 583.180 1049.200 ;
        RECT 582.920 765.040 583.180 765.300 ;
        RECT 605.920 765.040 606.180 765.300 ;
      LAYER met2 ;
        RECT 16.660 1049.085 16.920 1049.230 ;
        RECT 16.650 1048.715 16.930 1049.085 ;
        RECT 582.920 1048.910 583.180 1049.230 ;
        RECT 582.980 765.330 583.120 1048.910 ;
        RECT 582.920 765.010 583.180 765.330 ;
        RECT 605.920 765.010 606.180 765.330 ;
        RECT 605.980 749.770 606.120 765.010 ;
        RECT 606.630 749.770 606.910 750.000 ;
        RECT 605.980 749.630 606.910 749.770 ;
        RECT 606.630 746.000 606.910 749.630 ;
      LAYER via2 ;
        RECT 16.650 1048.760 16.930 1049.040 ;
      LAYER met3 ;
        RECT -4.800 1049.050 2.400 1049.500 ;
        RECT 16.625 1049.050 16.955 1049.065 ;
        RECT -4.800 1048.750 16.955 1049.050 ;
        RECT -4.800 1048.300 2.400 1048.750 ;
        RECT 16.625 1048.735 16.955 1048.750 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 793.800 16.030 793.860 ;
        RECT 582.430 793.800 582.750 793.860 ;
        RECT 15.710 793.660 582.750 793.800 ;
        RECT 15.710 793.600 16.030 793.660 ;
        RECT 582.430 793.600 582.750 793.660 ;
        RECT 582.430 764.900 582.750 764.960 ;
        RECT 610.030 764.900 610.350 764.960 ;
        RECT 582.430 764.760 610.350 764.900 ;
        RECT 582.430 764.700 582.750 764.760 ;
        RECT 610.030 764.700 610.350 764.760 ;
      LAYER via ;
        RECT 15.740 793.600 16.000 793.860 ;
        RECT 582.460 793.600 582.720 793.860 ;
        RECT 582.460 764.700 582.720 764.960 ;
        RECT 610.060 764.700 610.320 764.960 ;
      LAYER met2 ;
        RECT 15.730 797.795 16.010 798.165 ;
        RECT 15.800 793.890 15.940 797.795 ;
        RECT 15.740 793.570 16.000 793.890 ;
        RECT 582.460 793.570 582.720 793.890 ;
        RECT 582.520 764.990 582.660 793.570 ;
        RECT 582.460 764.670 582.720 764.990 ;
        RECT 610.060 764.670 610.320 764.990 ;
        RECT 610.120 749.770 610.260 764.670 ;
        RECT 610.770 749.770 611.050 750.000 ;
        RECT 610.120 749.630 611.050 749.770 ;
        RECT 610.770 746.000 611.050 749.630 ;
      LAYER via2 ;
        RECT 15.730 797.840 16.010 798.120 ;
      LAYER met3 ;
        RECT -4.800 798.130 2.400 798.580 ;
        RECT 15.705 798.130 16.035 798.145 ;
        RECT -4.800 797.830 16.035 798.130 ;
        RECT -4.800 797.380 2.400 797.830 ;
        RECT 15.705 797.815 16.035 797.830 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 763.540 614.490 763.600 ;
        RECT 590.800 763.400 614.490 763.540 ;
        RECT 23.990 762.180 24.310 762.240 ;
        RECT 590.800 762.180 590.940 763.400 ;
        RECT 614.170 763.340 614.490 763.400 ;
        RECT 23.990 762.040 590.940 762.180 ;
        RECT 23.990 761.980 24.310 762.040 ;
        RECT 13.870 550.700 14.190 550.760 ;
        RECT 23.990 550.700 24.310 550.760 ;
        RECT 13.870 550.560 24.310 550.700 ;
        RECT 13.870 550.500 14.190 550.560 ;
        RECT 23.990 550.500 24.310 550.560 ;
      LAYER via ;
        RECT 24.020 761.980 24.280 762.240 ;
        RECT 614.200 763.340 614.460 763.600 ;
        RECT 13.900 550.500 14.160 550.760 ;
        RECT 24.020 550.500 24.280 550.760 ;
      LAYER met2 ;
        RECT 614.200 763.310 614.460 763.630 ;
        RECT 24.020 761.950 24.280 762.270 ;
        RECT 24.080 550.790 24.220 761.950 ;
        RECT 614.260 749.770 614.400 763.310 ;
        RECT 614.910 749.770 615.190 750.000 ;
        RECT 614.260 749.630 615.190 749.770 ;
        RECT 614.910 746.000 615.190 749.630 ;
        RECT 13.900 550.470 14.160 550.790 ;
        RECT 24.020 550.470 24.280 550.790 ;
        RECT 13.960 547.245 14.100 550.470 ;
        RECT 13.890 546.875 14.170 547.245 ;
      LAYER via2 ;
        RECT 13.890 546.920 14.170 547.200 ;
      LAYER met3 ;
        RECT -4.800 547.210 2.400 547.660 ;
        RECT 13.865 547.210 14.195 547.225 ;
        RECT -4.800 546.910 14.195 547.210 ;
        RECT -4.800 546.460 2.400 546.910 ;
        RECT 13.865 546.895 14.195 546.910 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 753.340 18.790 753.400 ;
        RECT 618.310 753.340 618.630 753.400 ;
        RECT 18.470 753.200 618.630 753.340 ;
        RECT 18.470 753.140 18.790 753.200 ;
        RECT 618.310 753.140 618.630 753.200 ;
      LAYER via ;
        RECT 18.500 753.140 18.760 753.400 ;
        RECT 618.340 753.140 618.600 753.400 ;
      LAYER met2 ;
        RECT 18.500 753.110 18.760 753.430 ;
        RECT 618.340 753.110 618.600 753.430 ;
        RECT 18.560 296.325 18.700 753.110 ;
        RECT 618.400 749.770 618.540 753.110 ;
        RECT 619.050 749.770 619.330 750.000 ;
        RECT 618.400 749.630 619.330 749.770 ;
        RECT 619.050 746.000 619.330 749.630 ;
        RECT 18.490 295.955 18.770 296.325 ;
      LAYER via2 ;
        RECT 18.490 296.000 18.770 296.280 ;
      LAYER met3 ;
        RECT -4.800 296.290 2.400 296.740 ;
        RECT 18.465 296.290 18.795 296.305 ;
        RECT -4.800 295.990 18.795 296.290 ;
        RECT -4.800 295.540 2.400 295.990 ;
        RECT 18.465 295.975 18.795 295.990 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 752.660 16.490 752.720 ;
        RECT 622.450 752.660 622.770 752.720 ;
        RECT 16.170 752.520 622.770 752.660 ;
        RECT 16.170 752.460 16.490 752.520 ;
        RECT 622.450 752.460 622.770 752.520 ;
      LAYER via ;
        RECT 16.200 752.460 16.460 752.720 ;
        RECT 622.480 752.460 622.740 752.720 ;
      LAYER met2 ;
        RECT 16.200 752.430 16.460 752.750 ;
        RECT 622.480 752.430 622.740 752.750 ;
        RECT 16.260 711.010 16.400 752.430 ;
        RECT 622.540 749.770 622.680 752.430 ;
        RECT 623.190 749.770 623.470 750.000 ;
        RECT 622.540 749.630 623.470 749.770 ;
        RECT 623.190 746.000 623.470 749.630 ;
        RECT 16.260 710.870 17.320 711.010 ;
        RECT 17.180 45.405 17.320 710.870 ;
        RECT 17.110 45.035 17.390 45.405 ;
      LAYER via2 ;
        RECT 17.110 45.080 17.390 45.360 ;
      LAYER met3 ;
        RECT -4.800 45.370 2.400 45.820 ;
        RECT 17.085 45.370 17.415 45.385 ;
        RECT -4.800 45.070 17.415 45.370 ;
        RECT -4.800 44.620 2.400 45.070 ;
        RECT 17.085 45.055 17.415 45.070 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 897.160 443.370 897.220 ;
        RECT 2900.830 897.160 2901.150 897.220 ;
        RECT 443.050 897.020 2901.150 897.160 ;
        RECT 443.050 896.960 443.370 897.020 ;
        RECT 2900.830 896.960 2901.150 897.020 ;
      LAYER via ;
        RECT 443.080 896.960 443.340 897.220 ;
        RECT 2900.860 896.960 2901.120 897.220 ;
      LAYER met2 ;
        RECT 2900.850 899.115 2901.130 899.485 ;
        RECT 2900.920 897.250 2901.060 899.115 ;
        RECT 443.080 896.930 443.340 897.250 ;
        RECT 2900.860 896.930 2901.120 897.250 ;
        RECT 443.140 749.770 443.280 896.930 ;
        RECT 443.790 749.770 444.070 750.000 ;
        RECT 443.140 749.630 444.070 749.770 ;
        RECT 443.790 746.000 444.070 749.630 ;
      LAYER via2 ;
        RECT 2900.850 899.160 2901.130 899.440 ;
      LAYER met3 ;
        RECT 2900.825 899.450 2901.155 899.465 ;
        RECT 2917.600 899.450 2924.800 899.900 ;
        RECT 2900.825 899.150 2924.800 899.450 ;
        RECT 2900.825 899.135 2901.155 899.150 ;
        RECT 2917.600 898.700 2924.800 899.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 1131.760 449.350 1131.820 ;
        RECT 2900.830 1131.760 2901.150 1131.820 ;
        RECT 449.030 1131.620 2901.150 1131.760 ;
        RECT 449.030 1131.560 449.350 1131.620 ;
        RECT 2900.830 1131.560 2901.150 1131.620 ;
      LAYER via ;
        RECT 449.060 1131.560 449.320 1131.820 ;
        RECT 2900.860 1131.560 2901.120 1131.820 ;
      LAYER met2 ;
        RECT 2900.850 1133.715 2901.130 1134.085 ;
        RECT 2900.920 1131.850 2901.060 1133.715 ;
        RECT 449.060 1131.530 449.320 1131.850 ;
        RECT 2900.860 1131.530 2901.120 1131.850 ;
        RECT 449.120 751.130 449.260 1131.530 ;
        RECT 449.120 750.990 449.490 751.130 ;
        RECT 449.350 750.000 449.490 750.990 ;
        RECT 449.310 746.000 449.590 750.000 ;
      LAYER via2 ;
        RECT 2900.850 1133.760 2901.130 1134.040 ;
      LAYER met3 ;
        RECT 2900.825 1134.050 2901.155 1134.065 ;
        RECT 2917.600 1134.050 2924.800 1134.500 ;
        RECT 2900.825 1133.750 2924.800 1134.050 ;
        RECT 2900.825 1133.735 2901.155 1133.750 ;
        RECT 2917.600 1133.300 2924.800 1133.750 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 1366.360 448.890 1366.420 ;
        RECT 2900.830 1366.360 2901.150 1366.420 ;
        RECT 448.570 1366.220 2901.150 1366.360 ;
        RECT 448.570 1366.160 448.890 1366.220 ;
        RECT 2900.830 1366.160 2901.150 1366.220 ;
        RECT 448.570 766.260 448.890 766.320 ;
        RECT 454.090 766.260 454.410 766.320 ;
        RECT 448.570 766.120 454.410 766.260 ;
        RECT 448.570 766.060 448.890 766.120 ;
        RECT 454.090 766.060 454.410 766.120 ;
      LAYER via ;
        RECT 448.600 1366.160 448.860 1366.420 ;
        RECT 2900.860 1366.160 2901.120 1366.420 ;
        RECT 448.600 766.060 448.860 766.320 ;
        RECT 454.120 766.060 454.380 766.320 ;
      LAYER met2 ;
        RECT 2900.850 1368.315 2901.130 1368.685 ;
        RECT 2900.920 1366.450 2901.060 1368.315 ;
        RECT 448.600 1366.130 448.860 1366.450 ;
        RECT 2900.860 1366.130 2901.120 1366.450 ;
        RECT 448.660 766.350 448.800 1366.130 ;
        RECT 448.600 766.030 448.860 766.350 ;
        RECT 454.120 766.030 454.380 766.350 ;
        RECT 454.180 749.770 454.320 766.030 ;
        RECT 454.830 749.770 455.110 750.000 ;
        RECT 454.180 749.630 455.110 749.770 ;
        RECT 454.830 746.000 455.110 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1368.360 2901.130 1368.640 ;
      LAYER met3 ;
        RECT 2900.825 1368.650 2901.155 1368.665 ;
        RECT 2917.600 1368.650 2924.800 1369.100 ;
        RECT 2900.825 1368.350 2924.800 1368.650 ;
        RECT 2900.825 1368.335 2901.155 1368.350 ;
        RECT 2917.600 1367.900 2924.800 1368.350 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 1600.960 455.790 1601.020 ;
        RECT 2900.830 1600.960 2901.150 1601.020 ;
        RECT 455.470 1600.820 2901.150 1600.960 ;
        RECT 455.470 1600.760 455.790 1600.820 ;
        RECT 2900.830 1600.760 2901.150 1600.820 ;
        RECT 455.470 766.260 455.790 766.320 ;
        RECT 459.610 766.260 459.930 766.320 ;
        RECT 455.470 766.120 459.930 766.260 ;
        RECT 455.470 766.060 455.790 766.120 ;
        RECT 459.610 766.060 459.930 766.120 ;
      LAYER via ;
        RECT 455.500 1600.760 455.760 1601.020 ;
        RECT 2900.860 1600.760 2901.120 1601.020 ;
        RECT 455.500 766.060 455.760 766.320 ;
        RECT 459.640 766.060 459.900 766.320 ;
      LAYER met2 ;
        RECT 2900.850 1602.915 2901.130 1603.285 ;
        RECT 2900.920 1601.050 2901.060 1602.915 ;
        RECT 455.500 1600.730 455.760 1601.050 ;
        RECT 2900.860 1600.730 2901.120 1601.050 ;
        RECT 455.560 766.350 455.700 1600.730 ;
        RECT 455.500 766.030 455.760 766.350 ;
        RECT 459.640 766.030 459.900 766.350 ;
        RECT 459.700 749.770 459.840 766.030 ;
        RECT 460.350 749.770 460.630 750.000 ;
        RECT 459.700 749.630 460.630 749.770 ;
        RECT 460.350 746.000 460.630 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1602.960 2901.130 1603.240 ;
      LAYER met3 ;
        RECT 2900.825 1603.250 2901.155 1603.265 ;
        RECT 2917.600 1603.250 2924.800 1603.700 ;
        RECT 2900.825 1602.950 2924.800 1603.250 ;
        RECT 2900.825 1602.935 2901.155 1602.950 ;
        RECT 2917.600 1602.500 2924.800 1602.950 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 1835.560 462.690 1835.620 ;
        RECT 2900.830 1835.560 2901.150 1835.620 ;
        RECT 462.370 1835.420 2901.150 1835.560 ;
        RECT 462.370 1835.360 462.690 1835.420 ;
        RECT 2900.830 1835.360 2901.150 1835.420 ;
        RECT 462.370 766.600 462.690 766.660 ;
        RECT 465.130 766.600 465.450 766.660 ;
        RECT 462.370 766.460 465.450 766.600 ;
        RECT 462.370 766.400 462.690 766.460 ;
        RECT 465.130 766.400 465.450 766.460 ;
      LAYER via ;
        RECT 462.400 1835.360 462.660 1835.620 ;
        RECT 2900.860 1835.360 2901.120 1835.620 ;
        RECT 462.400 766.400 462.660 766.660 ;
        RECT 465.160 766.400 465.420 766.660 ;
      LAYER met2 ;
        RECT 2900.850 1837.515 2901.130 1837.885 ;
        RECT 2900.920 1835.650 2901.060 1837.515 ;
        RECT 462.400 1835.330 462.660 1835.650 ;
        RECT 2900.860 1835.330 2901.120 1835.650 ;
        RECT 462.460 766.690 462.600 1835.330 ;
        RECT 462.400 766.370 462.660 766.690 ;
        RECT 465.160 766.370 465.420 766.690 ;
        RECT 465.220 749.770 465.360 766.370 ;
        RECT 465.870 749.770 466.150 750.000 ;
        RECT 465.220 749.630 466.150 749.770 ;
        RECT 465.870 746.000 466.150 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1837.560 2901.130 1837.840 ;
      LAYER met3 ;
        RECT 2900.825 1837.850 2901.155 1837.865 ;
        RECT 2917.600 1837.850 2924.800 1838.300 ;
        RECT 2900.825 1837.550 2924.800 1837.850 ;
        RECT 2900.825 1837.535 2901.155 1837.550 ;
        RECT 2917.600 1837.100 2924.800 1837.550 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.650 2070.160 470.970 2070.220 ;
        RECT 2900.830 2070.160 2901.150 2070.220 ;
        RECT 470.650 2070.020 2901.150 2070.160 ;
        RECT 470.650 2069.960 470.970 2070.020 ;
        RECT 2900.830 2069.960 2901.150 2070.020 ;
      LAYER via ;
        RECT 470.680 2069.960 470.940 2070.220 ;
        RECT 2900.860 2069.960 2901.120 2070.220 ;
      LAYER met2 ;
        RECT 2900.850 2072.115 2901.130 2072.485 ;
        RECT 2900.920 2070.250 2901.060 2072.115 ;
        RECT 470.680 2069.930 470.940 2070.250 ;
        RECT 2900.860 2069.930 2901.120 2070.250 ;
        RECT 470.740 749.770 470.880 2069.930 ;
        RECT 471.390 749.770 471.670 750.000 ;
        RECT 470.740 749.630 471.670 749.770 ;
        RECT 471.390 746.000 471.670 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2072.160 2901.130 2072.440 ;
      LAYER met3 ;
        RECT 2900.825 2072.450 2901.155 2072.465 ;
        RECT 2917.600 2072.450 2924.800 2072.900 ;
        RECT 2900.825 2072.150 2924.800 2072.450 ;
        RECT 2900.825 2072.135 2901.155 2072.150 ;
        RECT 2917.600 2071.700 2924.800 2072.150 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.630 2304.760 476.950 2304.820 ;
        RECT 2900.830 2304.760 2901.150 2304.820 ;
        RECT 476.630 2304.620 2901.150 2304.760 ;
        RECT 476.630 2304.560 476.950 2304.620 ;
        RECT 2900.830 2304.560 2901.150 2304.620 ;
      LAYER via ;
        RECT 476.660 2304.560 476.920 2304.820 ;
        RECT 2900.860 2304.560 2901.120 2304.820 ;
      LAYER met2 ;
        RECT 2900.850 2306.715 2901.130 2307.085 ;
        RECT 2900.920 2304.850 2901.060 2306.715 ;
        RECT 476.660 2304.530 476.920 2304.850 ;
        RECT 2900.860 2304.530 2901.120 2304.850 ;
        RECT 476.720 751.130 476.860 2304.530 ;
        RECT 476.720 750.990 477.090 751.130 ;
        RECT 476.950 750.000 477.090 750.990 ;
        RECT 476.910 746.000 477.190 750.000 ;
      LAYER via2 ;
        RECT 2900.850 2306.760 2901.130 2307.040 ;
      LAYER met3 ;
        RECT 2900.825 2307.050 2901.155 2307.065 ;
        RECT 2917.600 2307.050 2924.800 2307.500 ;
        RECT 2900.825 2306.750 2924.800 2307.050 ;
        RECT 2900.825 2306.735 2901.155 2306.750 ;
        RECT 2917.600 2306.300 2924.800 2306.750 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.250 760.140 429.570 760.200 ;
        RECT 476.170 760.140 476.490 760.200 ;
        RECT 429.250 760.000 476.490 760.140 ;
        RECT 429.250 759.940 429.570 760.000 ;
        RECT 476.170 759.940 476.490 760.000 ;
        RECT 476.170 755.380 476.490 755.440 ;
        RECT 2901.750 755.380 2902.070 755.440 ;
        RECT 476.170 755.240 2902.070 755.380 ;
        RECT 476.170 755.180 476.490 755.240 ;
        RECT 2901.750 755.180 2902.070 755.240 ;
      LAYER via ;
        RECT 429.280 759.940 429.540 760.200 ;
        RECT 476.200 759.940 476.460 760.200 ;
        RECT 476.200 755.180 476.460 755.440 ;
        RECT 2901.780 755.180 2902.040 755.440 ;
      LAYER met2 ;
        RECT 429.280 759.910 429.540 760.230 ;
        RECT 476.200 759.910 476.460 760.230 ;
        RECT 428.610 749.770 428.890 750.000 ;
        RECT 429.340 749.770 429.480 759.910 ;
        RECT 476.260 755.470 476.400 759.910 ;
        RECT 476.200 755.150 476.460 755.470 ;
        RECT 2901.780 755.150 2902.040 755.470 ;
        RECT 428.610 749.630 429.480 749.770 ;
        RECT 428.610 746.000 428.890 749.630 ;
        RECT 2901.840 117.485 2901.980 755.150 ;
        RECT 2901.770 117.115 2902.050 117.485 ;
      LAYER via2 ;
        RECT 2901.770 117.160 2902.050 117.440 ;
      LAYER met3 ;
        RECT 2901.745 117.450 2902.075 117.465 ;
        RECT 2917.600 117.450 2924.800 117.900 ;
        RECT 2901.745 117.150 2924.800 117.450 ;
        RECT 2901.745 117.135 2902.075 117.150 ;
        RECT 2917.600 116.700 2924.800 117.150 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 2463.540 483.850 2463.600 ;
        RECT 2900.830 2463.540 2901.150 2463.600 ;
        RECT 483.530 2463.400 2901.150 2463.540 ;
        RECT 483.530 2463.340 483.850 2463.400 ;
        RECT 2900.830 2463.340 2901.150 2463.400 ;
      LAYER via ;
        RECT 483.560 2463.340 483.820 2463.600 ;
        RECT 2900.860 2463.340 2901.120 2463.600 ;
      LAYER met2 ;
        RECT 483.560 2463.310 483.820 2463.630 ;
        RECT 2900.860 2463.485 2901.120 2463.630 ;
        RECT 483.620 751.130 483.760 2463.310 ;
        RECT 2900.850 2463.115 2901.130 2463.485 ;
        RECT 483.620 750.990 483.990 751.130 ;
        RECT 483.850 750.000 483.990 750.990 ;
        RECT 483.810 746.000 484.090 750.000 ;
      LAYER via2 ;
        RECT 2900.850 2463.160 2901.130 2463.440 ;
      LAYER met3 ;
        RECT 2900.825 2463.450 2901.155 2463.465 ;
        RECT 2917.600 2463.450 2924.800 2463.900 ;
        RECT 2900.825 2463.150 2924.800 2463.450 ;
        RECT 2900.825 2463.135 2901.155 2463.150 ;
        RECT 2917.600 2462.700 2924.800 2463.150 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.450 2698.140 484.770 2698.200 ;
        RECT 2900.830 2698.140 2901.150 2698.200 ;
        RECT 484.450 2698.000 2901.150 2698.140 ;
        RECT 484.450 2697.940 484.770 2698.000 ;
        RECT 2900.830 2697.940 2901.150 2698.000 ;
        RECT 484.450 766.600 484.770 766.660 ;
        RECT 488.590 766.600 488.910 766.660 ;
        RECT 484.450 766.460 488.910 766.600 ;
        RECT 484.450 766.400 484.770 766.460 ;
        RECT 488.590 766.400 488.910 766.460 ;
      LAYER via ;
        RECT 484.480 2697.940 484.740 2698.200 ;
        RECT 2900.860 2697.940 2901.120 2698.200 ;
        RECT 484.480 766.400 484.740 766.660 ;
        RECT 488.620 766.400 488.880 766.660 ;
      LAYER met2 ;
        RECT 484.480 2697.910 484.740 2698.230 ;
        RECT 2900.860 2698.085 2901.120 2698.230 ;
        RECT 484.540 766.690 484.680 2697.910 ;
        RECT 2900.850 2697.715 2901.130 2698.085 ;
        RECT 484.480 766.370 484.740 766.690 ;
        RECT 488.620 766.370 488.880 766.690 ;
        RECT 488.680 749.770 488.820 766.370 ;
        RECT 489.330 749.770 489.610 750.000 ;
        RECT 488.680 749.630 489.610 749.770 ;
        RECT 489.330 746.000 489.610 749.630 ;
      LAYER via2 ;
        RECT 2900.850 2697.760 2901.130 2698.040 ;
      LAYER met3 ;
        RECT 2900.825 2698.050 2901.155 2698.065 ;
        RECT 2917.600 2698.050 2924.800 2698.500 ;
        RECT 2900.825 2697.750 2924.800 2698.050 ;
        RECT 2900.825 2697.735 2901.155 2697.750 ;
        RECT 2917.600 2697.300 2924.800 2697.750 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.350 2932.740 491.670 2932.800 ;
        RECT 2904.510 2932.740 2904.830 2932.800 ;
        RECT 491.350 2932.600 2904.830 2932.740 ;
        RECT 491.350 2932.540 491.670 2932.600 ;
        RECT 2904.510 2932.540 2904.830 2932.600 ;
        RECT 491.350 766.600 491.670 766.660 ;
        RECT 494.110 766.600 494.430 766.660 ;
        RECT 491.350 766.460 494.430 766.600 ;
        RECT 491.350 766.400 491.670 766.460 ;
        RECT 494.110 766.400 494.430 766.460 ;
      LAYER via ;
        RECT 491.380 2932.540 491.640 2932.800 ;
        RECT 2904.540 2932.540 2904.800 2932.800 ;
        RECT 491.380 766.400 491.640 766.660 ;
        RECT 494.140 766.400 494.400 766.660 ;
      LAYER met2 ;
        RECT 491.380 2932.510 491.640 2932.830 ;
        RECT 2904.540 2932.685 2904.800 2932.830 ;
        RECT 491.440 766.690 491.580 2932.510 ;
        RECT 2904.530 2932.315 2904.810 2932.685 ;
        RECT 491.380 766.370 491.640 766.690 ;
        RECT 494.140 766.370 494.400 766.690 ;
        RECT 494.200 749.770 494.340 766.370 ;
        RECT 494.850 749.770 495.130 750.000 ;
        RECT 494.200 749.630 495.130 749.770 ;
        RECT 494.850 746.000 495.130 749.630 ;
      LAYER via2 ;
        RECT 2904.530 2932.360 2904.810 2932.640 ;
      LAYER met3 ;
        RECT 2904.505 2932.650 2904.835 2932.665 ;
        RECT 2917.600 2932.650 2924.800 2933.100 ;
        RECT 2904.505 2932.335 2905.050 2932.650 ;
        RECT 2904.750 2931.970 2905.050 2932.335 ;
        RECT 2914.870 2932.350 2924.800 2932.650 ;
        RECT 2914.870 2931.970 2915.170 2932.350 ;
        RECT 2904.750 2931.670 2915.170 2931.970 ;
        RECT 2917.600 2931.900 2924.800 2932.350 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 499.630 3167.340 499.950 3167.400 ;
        RECT 2900.830 3167.340 2901.150 3167.400 ;
        RECT 499.630 3167.200 2901.150 3167.340 ;
        RECT 499.630 3167.140 499.950 3167.200 ;
        RECT 2900.830 3167.140 2901.150 3167.200 ;
      LAYER via ;
        RECT 499.660 3167.140 499.920 3167.400 ;
        RECT 2900.860 3167.140 2901.120 3167.400 ;
      LAYER met2 ;
        RECT 499.660 3167.110 499.920 3167.430 ;
        RECT 2900.860 3167.285 2901.120 3167.430 ;
        RECT 499.720 749.770 499.860 3167.110 ;
        RECT 2900.850 3166.915 2901.130 3167.285 ;
        RECT 500.370 749.770 500.650 750.000 ;
        RECT 499.720 749.630 500.650 749.770 ;
        RECT 500.370 746.000 500.650 749.630 ;
      LAYER via2 ;
        RECT 2900.850 3166.960 2901.130 3167.240 ;
      LAYER met3 ;
        RECT 2900.825 3167.250 2901.155 3167.265 ;
        RECT 2917.600 3167.250 2924.800 3167.700 ;
        RECT 2900.825 3166.950 2924.800 3167.250 ;
        RECT 2900.825 3166.935 2901.155 3166.950 ;
        RECT 2917.600 3166.500 2924.800 3166.950 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 505.150 3401.940 505.470 3402.000 ;
        RECT 2900.830 3401.940 2901.150 3402.000 ;
        RECT 505.150 3401.800 2901.150 3401.940 ;
        RECT 505.150 3401.740 505.470 3401.800 ;
        RECT 2900.830 3401.740 2901.150 3401.800 ;
      LAYER via ;
        RECT 505.180 3401.740 505.440 3402.000 ;
        RECT 2900.860 3401.740 2901.120 3402.000 ;
      LAYER met2 ;
        RECT 505.180 3401.710 505.440 3402.030 ;
        RECT 2900.860 3401.885 2901.120 3402.030 ;
        RECT 505.240 749.770 505.380 3401.710 ;
        RECT 2900.850 3401.515 2901.130 3401.885 ;
        RECT 505.890 749.770 506.170 750.000 ;
        RECT 505.240 749.630 506.170 749.770 ;
        RECT 505.890 746.000 506.170 749.630 ;
      LAYER via2 ;
        RECT 2900.850 3401.560 2901.130 3401.840 ;
      LAYER met3 ;
        RECT 2900.825 3401.850 2901.155 3401.865 ;
        RECT 2917.600 3401.850 2924.800 3402.300 ;
        RECT 2900.825 3401.550 2924.800 3401.850 ;
        RECT 2900.825 3401.535 2901.155 3401.550 ;
        RECT 2917.600 3401.100 2924.800 3401.550 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 3501.560 511.450 3501.620 ;
        RECT 2756.850 3501.560 2757.170 3501.620 ;
        RECT 511.130 3501.420 2757.170 3501.560 ;
        RECT 511.130 3501.360 511.450 3501.420 ;
        RECT 2756.850 3501.360 2757.170 3501.420 ;
      LAYER via ;
        RECT 511.160 3501.360 511.420 3501.620 ;
        RECT 2756.880 3501.360 2757.140 3501.620 ;
      LAYER met2 ;
        RECT 2756.730 3517.600 2757.290 3524.800 ;
        RECT 2756.940 3501.650 2757.080 3517.600 ;
        RECT 511.160 3501.330 511.420 3501.650 ;
        RECT 2756.880 3501.330 2757.140 3501.650 ;
        RECT 511.220 751.130 511.360 3501.330 ;
        RECT 511.220 750.990 511.590 751.130 ;
        RECT 511.450 750.000 511.590 750.990 ;
        RECT 511.410 746.000 511.690 750.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 3501.900 510.990 3501.960 ;
        RECT 2432.550 3501.900 2432.870 3501.960 ;
        RECT 510.670 3501.760 2432.870 3501.900 ;
        RECT 510.670 3501.700 510.990 3501.760 ;
        RECT 2432.550 3501.700 2432.870 3501.760 ;
        RECT 510.670 791.420 510.990 791.480 ;
        RECT 516.190 791.420 516.510 791.480 ;
        RECT 510.670 791.280 516.510 791.420 ;
        RECT 510.670 791.220 510.990 791.280 ;
        RECT 516.190 791.220 516.510 791.280 ;
      LAYER via ;
        RECT 510.700 3501.700 510.960 3501.960 ;
        RECT 2432.580 3501.700 2432.840 3501.960 ;
        RECT 510.700 791.220 510.960 791.480 ;
        RECT 516.220 791.220 516.480 791.480 ;
      LAYER met2 ;
        RECT 2432.430 3517.600 2432.990 3524.800 ;
        RECT 2432.640 3501.990 2432.780 3517.600 ;
        RECT 510.700 3501.670 510.960 3501.990 ;
        RECT 2432.580 3501.670 2432.840 3501.990 ;
        RECT 510.760 791.510 510.900 3501.670 ;
        RECT 510.700 791.190 510.960 791.510 ;
        RECT 516.220 791.190 516.480 791.510 ;
        RECT 516.280 749.770 516.420 791.190 ;
        RECT 516.930 749.770 517.210 750.000 ;
        RECT 516.280 749.630 517.210 749.770 ;
        RECT 516.930 746.000 517.210 749.630 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 3502.240 517.890 3502.300 ;
        RECT 2108.250 3502.240 2108.570 3502.300 ;
        RECT 517.570 3502.100 2108.570 3502.240 ;
        RECT 517.570 3502.040 517.890 3502.100 ;
        RECT 2108.250 3502.040 2108.570 3502.100 ;
      LAYER via ;
        RECT 517.600 3502.040 517.860 3502.300 ;
        RECT 2108.280 3502.040 2108.540 3502.300 ;
      LAYER met2 ;
        RECT 2108.130 3517.600 2108.690 3524.800 ;
        RECT 2108.340 3502.330 2108.480 3517.600 ;
        RECT 517.600 3502.010 517.860 3502.330 ;
        RECT 2108.280 3502.010 2108.540 3502.330 ;
        RECT 517.660 855.670 517.800 3502.010 ;
        RECT 517.660 855.530 521.940 855.670 ;
        RECT 521.800 749.770 521.940 855.530 ;
        RECT 522.450 749.770 522.730 750.000 ;
        RECT 521.800 749.630 522.730 749.770 ;
        RECT 522.450 746.000 522.730 749.630 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 783.260 527.550 783.320 ;
        RECT 1780.270 783.260 1780.590 783.320 ;
        RECT 527.230 783.120 1780.590 783.260 ;
        RECT 527.230 783.060 527.550 783.120 ;
        RECT 1780.270 783.060 1780.590 783.120 ;
      LAYER via ;
        RECT 527.260 783.060 527.520 783.320 ;
        RECT 1780.300 783.060 1780.560 783.320 ;
      LAYER met2 ;
        RECT 1780.360 3517.910 1783.260 3518.050 ;
        RECT 1780.360 783.350 1780.500 3517.910 ;
        RECT 1783.120 3517.370 1783.260 3517.910 ;
        RECT 1783.830 3517.600 1784.390 3524.800 ;
        RECT 1784.040 3517.370 1784.180 3517.600 ;
        RECT 1783.120 3517.230 1784.180 3517.370 ;
        RECT 527.260 783.030 527.520 783.350 ;
        RECT 1780.300 783.030 1780.560 783.350 ;
        RECT 527.320 749.770 527.460 783.030 ;
        RECT 527.970 749.770 528.250 750.000 ;
        RECT 527.320 749.630 528.250 749.770 ;
        RECT 527.970 746.000 528.250 749.630 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 3502.580 531.690 3502.640 ;
        RECT 1459.650 3502.580 1459.970 3502.640 ;
        RECT 531.370 3502.440 1459.970 3502.580 ;
        RECT 531.370 3502.380 531.690 3502.440 ;
        RECT 1459.650 3502.380 1459.970 3502.440 ;
      LAYER via ;
        RECT 531.400 3502.380 531.660 3502.640 ;
        RECT 1459.680 3502.380 1459.940 3502.640 ;
      LAYER met2 ;
        RECT 1459.530 3517.600 1460.090 3524.800 ;
        RECT 1459.740 3502.670 1459.880 3517.600 ;
        RECT 531.400 3502.350 531.660 3502.670 ;
        RECT 1459.680 3502.350 1459.940 3502.670 ;
        RECT 531.460 855.670 531.600 3502.350 ;
        RECT 531.460 855.530 532.980 855.670 ;
        RECT 532.840 749.770 532.980 855.530 ;
        RECT 533.490 749.770 533.770 750.000 ;
        RECT 532.840 749.630 533.770 749.770 ;
        RECT 533.490 746.000 533.770 749.630 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 680.410 358.600 680.730 358.660 ;
        RECT 2898.070 358.600 2898.390 358.660 ;
        RECT 680.410 358.460 2898.390 358.600 ;
        RECT 680.410 358.400 680.730 358.460 ;
        RECT 2898.070 358.400 2898.390 358.460 ;
      LAYER via ;
        RECT 680.440 358.400 680.700 358.660 ;
        RECT 2898.100 358.400 2898.360 358.660 ;
      LAYER met2 ;
        RECT 434.330 762.435 434.610 762.805 ;
        RECT 680.430 762.435 680.710 762.805 ;
        RECT 434.400 750.000 434.540 762.435 ;
        RECT 434.130 749.630 434.540 750.000 ;
        RECT 434.130 746.000 434.410 749.630 ;
        RECT 680.500 358.690 680.640 762.435 ;
        RECT 680.440 358.370 680.700 358.690 ;
        RECT 2898.100 358.370 2898.360 358.690 ;
        RECT 2898.160 352.085 2898.300 358.370 ;
        RECT 2898.090 351.715 2898.370 352.085 ;
      LAYER via2 ;
        RECT 434.330 762.480 434.610 762.760 ;
        RECT 680.430 762.480 680.710 762.760 ;
        RECT 2898.090 351.760 2898.370 352.040 ;
      LAYER met3 ;
        RECT 434.305 762.770 434.635 762.785 ;
        RECT 680.405 762.770 680.735 762.785 ;
        RECT 434.305 762.470 680.735 762.770 ;
        RECT 434.305 762.455 434.635 762.470 ;
        RECT 680.405 762.455 680.735 762.470 ;
        RECT 2898.065 352.050 2898.395 352.065 ;
        RECT 2917.600 352.050 2924.800 352.500 ;
        RECT 2898.065 351.750 2924.800 352.050 ;
        RECT 2898.065 351.735 2898.395 351.750 ;
        RECT 2917.600 351.300 2924.800 351.750 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 3502.920 539.050 3502.980 ;
        RECT 1135.350 3502.920 1135.670 3502.980 ;
        RECT 538.730 3502.780 1135.670 3502.920 ;
        RECT 538.730 3502.720 539.050 3502.780 ;
        RECT 1135.350 3502.720 1135.670 3502.780 ;
      LAYER via ;
        RECT 538.760 3502.720 539.020 3502.980 ;
        RECT 1135.380 3502.720 1135.640 3502.980 ;
      LAYER met2 ;
        RECT 1135.230 3517.600 1135.790 3524.800 ;
        RECT 1135.440 3503.010 1135.580 3517.600 ;
        RECT 538.760 3502.690 539.020 3503.010 ;
        RECT 1135.380 3502.690 1135.640 3503.010 ;
        RECT 538.820 751.130 538.960 3502.690 ;
        RECT 538.820 750.990 539.190 751.130 ;
        RECT 539.050 750.000 539.190 750.990 ;
        RECT 539.010 746.000 539.290 750.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 3503.600 538.590 3503.660 ;
        RECT 811.050 3503.600 811.370 3503.660 ;
        RECT 538.270 3503.460 811.370 3503.600 ;
        RECT 538.270 3503.400 538.590 3503.460 ;
        RECT 811.050 3503.400 811.370 3503.460 ;
        RECT 538.270 794.480 538.590 794.540 ;
        RECT 543.790 794.480 544.110 794.540 ;
        RECT 538.270 794.340 544.110 794.480 ;
        RECT 538.270 794.280 538.590 794.340 ;
        RECT 543.790 794.280 544.110 794.340 ;
      LAYER via ;
        RECT 538.300 3503.400 538.560 3503.660 ;
        RECT 811.080 3503.400 811.340 3503.660 ;
        RECT 538.300 794.280 538.560 794.540 ;
        RECT 543.820 794.280 544.080 794.540 ;
      LAYER met2 ;
        RECT 810.930 3517.600 811.490 3524.800 ;
        RECT 811.140 3503.690 811.280 3517.600 ;
        RECT 538.300 3503.370 538.560 3503.690 ;
        RECT 811.080 3503.370 811.340 3503.690 ;
        RECT 538.360 794.570 538.500 3503.370 ;
        RECT 538.300 794.250 538.560 794.570 ;
        RECT 543.820 794.250 544.080 794.570 ;
        RECT 543.880 749.770 544.020 794.250 ;
        RECT 544.530 749.770 544.810 750.000 ;
        RECT 543.880 749.630 544.810 749.770 ;
        RECT 544.530 746.000 544.810 749.630 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.750 3503.940 487.070 3504.000 ;
        RECT 545.170 3503.940 545.490 3504.000 ;
        RECT 486.750 3503.800 545.490 3503.940 ;
        RECT 486.750 3503.740 487.070 3503.800 ;
        RECT 545.170 3503.740 545.490 3503.800 ;
      LAYER via ;
        RECT 486.780 3503.740 487.040 3504.000 ;
        RECT 545.200 3503.740 545.460 3504.000 ;
      LAYER met2 ;
        RECT 486.630 3517.600 487.190 3524.800 ;
        RECT 486.840 3504.030 486.980 3517.600 ;
        RECT 486.780 3503.710 487.040 3504.030 ;
        RECT 545.200 3503.710 545.460 3504.030 ;
        RECT 545.260 855.670 545.400 3503.710 ;
        RECT 545.260 855.530 549.540 855.670 ;
        RECT 549.400 749.770 549.540 855.530 ;
        RECT 550.050 749.770 550.330 750.000 ;
        RECT 549.400 749.630 550.330 749.770 ;
        RECT 550.050 746.000 550.330 749.630 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 162.450 3503.260 162.770 3503.320 ;
        RECT 554.830 3503.260 555.150 3503.320 ;
        RECT 162.450 3503.120 555.150 3503.260 ;
        RECT 162.450 3503.060 162.770 3503.120 ;
        RECT 554.830 3503.060 555.150 3503.120 ;
      LAYER via ;
        RECT 162.480 3503.060 162.740 3503.320 ;
        RECT 554.860 3503.060 555.120 3503.320 ;
      LAYER met2 ;
        RECT 162.330 3517.600 162.890 3524.800 ;
        RECT 162.540 3503.350 162.680 3517.600 ;
        RECT 162.480 3503.030 162.740 3503.350 ;
        RECT 554.860 3503.030 555.120 3503.350 ;
        RECT 554.920 749.770 555.060 3503.030 ;
        RECT 555.570 749.770 555.850 750.000 ;
        RECT 554.920 749.630 555.850 749.770 ;
        RECT 555.570 746.000 555.850 749.630 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3388.000 17.410 3388.060 ;
        RECT 560.810 3388.000 561.130 3388.060 ;
        RECT 17.090 3387.860 561.130 3388.000 ;
        RECT 17.090 3387.800 17.410 3387.860 ;
        RECT 560.810 3387.800 561.130 3387.860 ;
      LAYER via ;
        RECT 17.120 3387.800 17.380 3388.060 ;
        RECT 560.840 3387.800 561.100 3388.060 ;
      LAYER met2 ;
        RECT 17.110 3390.635 17.390 3391.005 ;
        RECT 17.180 3388.090 17.320 3390.635 ;
        RECT 17.120 3387.770 17.380 3388.090 ;
        RECT 560.840 3387.770 561.100 3388.090 ;
        RECT 560.900 751.130 561.040 3387.770 ;
        RECT 560.900 750.990 561.270 751.130 ;
        RECT 561.130 750.000 561.270 750.990 ;
        RECT 561.090 746.000 561.370 750.000 ;
      LAYER via2 ;
        RECT 17.110 3390.680 17.390 3390.960 ;
      LAYER met3 ;
        RECT -4.800 3390.970 2.400 3391.420 ;
        RECT 17.085 3390.970 17.415 3390.985 ;
        RECT -4.800 3390.670 17.415 3390.970 ;
        RECT -4.800 3390.220 2.400 3390.670 ;
        RECT 17.085 3390.655 17.415 3390.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3139.800 17.410 3139.860 ;
        RECT 566.790 3139.800 567.110 3139.860 ;
        RECT 17.090 3139.660 567.110 3139.800 ;
        RECT 17.090 3139.600 17.410 3139.660 ;
        RECT 566.790 3139.600 567.110 3139.660 ;
      LAYER via ;
        RECT 17.120 3139.600 17.380 3139.860 ;
        RECT 566.820 3139.600 567.080 3139.860 ;
      LAYER met2 ;
        RECT 17.110 3139.715 17.390 3140.085 ;
        RECT 17.120 3139.570 17.380 3139.715 ;
        RECT 566.820 3139.570 567.080 3139.890 ;
        RECT 566.880 750.000 567.020 3139.570 ;
        RECT 566.610 749.630 567.020 750.000 ;
        RECT 566.610 746.000 566.890 749.630 ;
      LAYER via2 ;
        RECT 17.110 3139.760 17.390 3140.040 ;
      LAYER met3 ;
        RECT -4.800 3140.050 2.400 3140.500 ;
        RECT 17.085 3140.050 17.415 3140.065 ;
        RECT -4.800 3139.750 17.415 3140.050 ;
        RECT -4.800 3139.300 2.400 3139.750 ;
        RECT 17.085 3139.735 17.415 3139.750 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2884.460 15.570 2884.520 ;
        RECT 570.010 2884.460 570.330 2884.520 ;
        RECT 15.250 2884.320 570.330 2884.460 ;
        RECT 15.250 2884.260 15.570 2884.320 ;
        RECT 570.010 2884.260 570.330 2884.320 ;
      LAYER via ;
        RECT 15.280 2884.260 15.540 2884.520 ;
        RECT 570.040 2884.260 570.300 2884.520 ;
      LAYER met2 ;
        RECT 15.270 2888.795 15.550 2889.165 ;
        RECT 15.340 2884.550 15.480 2888.795 ;
        RECT 15.280 2884.230 15.540 2884.550 ;
        RECT 570.040 2884.230 570.300 2884.550 ;
        RECT 570.100 855.670 570.240 2884.230 ;
        RECT 570.100 855.530 571.620 855.670 ;
        RECT 571.480 749.770 571.620 855.530 ;
        RECT 572.130 749.770 572.410 750.000 ;
        RECT 571.480 749.630 572.410 749.770 ;
        RECT 572.130 746.000 572.410 749.630 ;
      LAYER via2 ;
        RECT 15.270 2888.840 15.550 2889.120 ;
      LAYER met3 ;
        RECT -4.800 2889.130 2.400 2889.580 ;
        RECT 15.245 2889.130 15.575 2889.145 ;
        RECT -4.800 2888.830 15.575 2889.130 ;
        RECT -4.800 2888.380 2.400 2888.830 ;
        RECT 15.245 2888.815 15.575 2888.830 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 2635.920 18.330 2635.980 ;
        RECT 575.530 2635.920 575.850 2635.980 ;
        RECT 18.010 2635.780 575.850 2635.920 ;
        RECT 18.010 2635.720 18.330 2635.780 ;
        RECT 575.530 2635.720 575.850 2635.780 ;
      LAYER via ;
        RECT 18.040 2635.720 18.300 2635.980 ;
        RECT 575.560 2635.720 575.820 2635.980 ;
      LAYER met2 ;
        RECT 18.030 2637.875 18.310 2638.245 ;
        RECT 18.100 2636.010 18.240 2637.875 ;
        RECT 18.040 2635.690 18.300 2636.010 ;
        RECT 575.560 2635.690 575.820 2636.010 ;
        RECT 575.620 759.070 575.760 2635.690 ;
        RECT 575.620 758.930 577.140 759.070 ;
        RECT 577.000 749.770 577.140 758.930 ;
        RECT 577.650 749.770 577.930 750.000 ;
        RECT 577.000 749.630 577.930 749.770 ;
        RECT 577.650 746.000 577.930 749.630 ;
      LAYER via2 ;
        RECT 18.030 2637.920 18.310 2638.200 ;
      LAYER met3 ;
        RECT -4.800 2638.210 2.400 2638.660 ;
        RECT 18.005 2638.210 18.335 2638.225 ;
        RECT -4.800 2637.910 18.335 2638.210 ;
        RECT -4.800 2637.460 2.400 2637.910 ;
        RECT 18.005 2637.895 18.335 2637.910 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2380.920 16.030 2380.980 ;
        RECT 583.810 2380.920 584.130 2380.980 ;
        RECT 15.710 2380.780 584.130 2380.920 ;
        RECT 15.710 2380.720 16.030 2380.780 ;
        RECT 583.810 2380.720 584.130 2380.780 ;
      LAYER via ;
        RECT 15.740 2380.720 16.000 2380.980 ;
        RECT 583.840 2380.720 584.100 2380.980 ;
      LAYER met2 ;
        RECT 15.730 2386.955 16.010 2387.325 ;
        RECT 15.800 2381.010 15.940 2386.955 ;
        RECT 15.740 2380.690 16.000 2381.010 ;
        RECT 583.840 2380.690 584.100 2381.010 ;
        RECT 583.170 749.770 583.450 750.000 ;
        RECT 583.900 749.770 584.040 2380.690 ;
        RECT 583.170 749.630 584.040 749.770 ;
        RECT 583.170 746.000 583.450 749.630 ;
      LAYER via2 ;
        RECT 15.730 2387.000 16.010 2387.280 ;
      LAYER met3 ;
        RECT -4.800 2387.290 2.400 2387.740 ;
        RECT 15.705 2387.290 16.035 2387.305 ;
        RECT -4.800 2386.990 16.035 2387.290 ;
        RECT -4.800 2386.540 2.400 2386.990 ;
        RECT 15.705 2386.975 16.035 2386.990 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2132.380 16.950 2132.440 ;
        RECT 587.950 2132.380 588.270 2132.440 ;
        RECT 16.630 2132.240 588.270 2132.380 ;
        RECT 16.630 2132.180 16.950 2132.240 ;
        RECT 587.950 2132.180 588.270 2132.240 ;
      LAYER via ;
        RECT 16.660 2132.180 16.920 2132.440 ;
        RECT 587.980 2132.180 588.240 2132.440 ;
      LAYER met2 ;
        RECT 16.650 2136.035 16.930 2136.405 ;
        RECT 16.720 2132.470 16.860 2136.035 ;
        RECT 16.660 2132.150 16.920 2132.470 ;
        RECT 587.980 2132.150 588.240 2132.470 ;
        RECT 588.040 749.770 588.180 2132.150 ;
        RECT 588.690 749.770 588.970 750.000 ;
        RECT 588.040 749.630 588.970 749.770 ;
        RECT 588.690 746.000 588.970 749.630 ;
      LAYER via2 ;
        RECT 16.650 2136.080 16.930 2136.360 ;
      LAYER met3 ;
        RECT -4.800 2136.370 2.400 2136.820 ;
        RECT 16.625 2136.370 16.955 2136.385 ;
        RECT -4.800 2136.070 16.955 2136.370 ;
        RECT -4.800 2135.620 2.400 2136.070 ;
        RECT 16.625 2136.055 16.955 2136.070 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 693.290 593.200 693.610 593.260 ;
        RECT 2900.830 593.200 2901.150 593.260 ;
        RECT 693.290 593.060 2901.150 593.200 ;
        RECT 693.290 593.000 693.610 593.060 ;
        RECT 2900.830 593.000 2901.150 593.060 ;
      LAYER via ;
        RECT 693.320 593.000 693.580 593.260 ;
        RECT 2900.860 593.000 2901.120 593.260 ;
      LAYER met2 ;
        RECT 440.310 761.755 440.590 762.125 ;
        RECT 693.310 761.755 693.590 762.125 ;
        RECT 439.650 749.770 439.930 750.000 ;
        RECT 440.380 749.770 440.520 761.755 ;
        RECT 439.650 749.630 440.520 749.770 ;
        RECT 439.650 746.000 439.930 749.630 ;
        RECT 693.380 593.290 693.520 761.755 ;
        RECT 693.320 592.970 693.580 593.290 ;
        RECT 2900.860 592.970 2901.120 593.290 ;
        RECT 2900.920 586.685 2901.060 592.970 ;
        RECT 2900.850 586.315 2901.130 586.685 ;
      LAYER via2 ;
        RECT 440.310 761.800 440.590 762.080 ;
        RECT 693.310 761.800 693.590 762.080 ;
        RECT 2900.850 586.360 2901.130 586.640 ;
      LAYER met3 ;
        RECT 440.285 762.090 440.615 762.105 ;
        RECT 693.285 762.090 693.615 762.105 ;
        RECT 440.285 761.790 693.615 762.090 ;
        RECT 440.285 761.775 440.615 761.790 ;
        RECT 693.285 761.775 693.615 761.790 ;
        RECT 2900.825 586.650 2901.155 586.665 ;
        RECT 2917.600 586.650 2924.800 587.100 ;
        RECT 2900.825 586.350 2924.800 586.650 ;
        RECT 2900.825 586.335 2901.155 586.350 ;
        RECT 2917.600 585.900 2924.800 586.350 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1883.840 16.950 1883.900 ;
        RECT 589.790 1883.840 590.110 1883.900 ;
        RECT 16.630 1883.700 590.110 1883.840 ;
        RECT 16.630 1883.640 16.950 1883.700 ;
        RECT 589.790 1883.640 590.110 1883.700 ;
        RECT 589.790 772.720 590.110 772.780 ;
        RECT 593.470 772.720 593.790 772.780 ;
        RECT 589.790 772.580 593.790 772.720 ;
        RECT 589.790 772.520 590.110 772.580 ;
        RECT 593.470 772.520 593.790 772.580 ;
      LAYER via ;
        RECT 16.660 1883.640 16.920 1883.900 ;
        RECT 589.820 1883.640 590.080 1883.900 ;
        RECT 589.820 772.520 590.080 772.780 ;
        RECT 593.500 772.520 593.760 772.780 ;
      LAYER met2 ;
        RECT 16.650 1885.115 16.930 1885.485 ;
        RECT 16.720 1883.930 16.860 1885.115 ;
        RECT 16.660 1883.610 16.920 1883.930 ;
        RECT 589.820 1883.610 590.080 1883.930 ;
        RECT 589.880 772.810 590.020 1883.610 ;
        RECT 589.820 772.490 590.080 772.810 ;
        RECT 593.500 772.490 593.760 772.810 ;
        RECT 593.560 749.770 593.700 772.490 ;
        RECT 594.210 749.770 594.490 750.000 ;
        RECT 593.560 749.630 594.490 749.770 ;
        RECT 594.210 746.000 594.490 749.630 ;
      LAYER via2 ;
        RECT 16.650 1885.160 16.930 1885.440 ;
      LAYER met3 ;
        RECT -4.800 1885.450 2.400 1885.900 ;
        RECT 16.625 1885.450 16.955 1885.465 ;
        RECT -4.800 1885.150 16.955 1885.450 ;
        RECT -4.800 1884.700 2.400 1885.150 ;
        RECT 16.625 1885.135 16.955 1885.150 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1628.500 16.950 1628.560 ;
        RECT 590.250 1628.500 590.570 1628.560 ;
        RECT 16.630 1628.360 590.570 1628.500 ;
        RECT 16.630 1628.300 16.950 1628.360 ;
        RECT 590.250 1628.300 590.570 1628.360 ;
        RECT 590.250 779.520 590.570 779.580 ;
        RECT 598.990 779.520 599.310 779.580 ;
        RECT 590.250 779.380 599.310 779.520 ;
        RECT 590.250 779.320 590.570 779.380 ;
        RECT 598.990 779.320 599.310 779.380 ;
      LAYER via ;
        RECT 16.660 1628.300 16.920 1628.560 ;
        RECT 590.280 1628.300 590.540 1628.560 ;
        RECT 590.280 779.320 590.540 779.580 ;
        RECT 599.020 779.320 599.280 779.580 ;
      LAYER met2 ;
        RECT 16.650 1634.195 16.930 1634.565 ;
        RECT 16.720 1628.590 16.860 1634.195 ;
        RECT 16.660 1628.270 16.920 1628.590 ;
        RECT 590.280 1628.270 590.540 1628.590 ;
        RECT 590.340 779.610 590.480 1628.270 ;
        RECT 590.280 779.290 590.540 779.610 ;
        RECT 599.020 779.290 599.280 779.610 ;
        RECT 599.080 749.770 599.220 779.290 ;
        RECT 599.730 749.770 600.010 750.000 ;
        RECT 599.080 749.630 600.010 749.770 ;
        RECT 599.730 746.000 600.010 749.630 ;
      LAYER via2 ;
        RECT 16.650 1634.240 16.930 1634.520 ;
      LAYER met3 ;
        RECT -4.800 1634.530 2.400 1634.980 ;
        RECT 16.625 1634.530 16.955 1634.545 ;
        RECT -4.800 1634.230 16.955 1634.530 ;
        RECT -4.800 1633.780 2.400 1634.230 ;
        RECT 16.625 1634.215 16.955 1634.230 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1380.300 16.950 1380.360 ;
        RECT 603.590 1380.300 603.910 1380.360 ;
        RECT 16.630 1380.160 603.910 1380.300 ;
        RECT 16.630 1380.100 16.950 1380.160 ;
        RECT 603.590 1380.100 603.910 1380.160 ;
      LAYER via ;
        RECT 16.660 1380.100 16.920 1380.360 ;
        RECT 603.620 1380.100 603.880 1380.360 ;
      LAYER met2 ;
        RECT 16.650 1383.275 16.930 1383.645 ;
        RECT 16.720 1380.390 16.860 1383.275 ;
        RECT 16.660 1380.070 16.920 1380.390 ;
        RECT 603.620 1380.070 603.880 1380.390 ;
        RECT 603.680 751.130 603.820 1380.070 ;
        RECT 603.680 750.990 604.050 751.130 ;
        RECT 603.910 750.000 604.050 750.990 ;
        RECT 603.870 746.000 604.150 750.000 ;
      LAYER via2 ;
        RECT 16.650 1383.320 16.930 1383.600 ;
      LAYER met3 ;
        RECT -4.800 1383.610 2.400 1384.060 ;
        RECT 16.625 1383.610 16.955 1383.625 ;
        RECT -4.800 1383.310 16.955 1383.610 ;
        RECT -4.800 1382.860 2.400 1383.310 ;
        RECT 16.625 1383.295 16.955 1383.310 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1132.100 16.950 1132.160 ;
        RECT 590.710 1132.100 591.030 1132.160 ;
        RECT 16.630 1131.960 591.030 1132.100 ;
        RECT 16.630 1131.900 16.950 1131.960 ;
        RECT 590.710 1131.900 591.030 1131.960 ;
        RECT 590.710 765.920 591.030 765.980 ;
        RECT 607.270 765.920 607.590 765.980 ;
        RECT 590.710 765.780 607.590 765.920 ;
        RECT 590.710 765.720 591.030 765.780 ;
        RECT 607.270 765.720 607.590 765.780 ;
      LAYER via ;
        RECT 16.660 1131.900 16.920 1132.160 ;
        RECT 590.740 1131.900 591.000 1132.160 ;
        RECT 590.740 765.720 591.000 765.980 ;
        RECT 607.300 765.720 607.560 765.980 ;
      LAYER met2 ;
        RECT 16.650 1132.355 16.930 1132.725 ;
        RECT 16.720 1132.190 16.860 1132.355 ;
        RECT 16.660 1131.870 16.920 1132.190 ;
        RECT 590.740 1131.870 591.000 1132.190 ;
        RECT 590.800 766.010 590.940 1131.870 ;
        RECT 590.740 765.690 591.000 766.010 ;
        RECT 607.300 765.690 607.560 766.010 ;
        RECT 607.360 749.770 607.500 765.690 ;
        RECT 608.010 749.770 608.290 750.000 ;
        RECT 607.360 749.630 608.290 749.770 ;
        RECT 608.010 746.000 608.290 749.630 ;
      LAYER via2 ;
        RECT 16.650 1132.400 16.930 1132.680 ;
      LAYER met3 ;
        RECT -4.800 1132.690 2.400 1133.140 ;
        RECT 16.625 1132.690 16.955 1132.705 ;
        RECT -4.800 1132.390 16.955 1132.690 ;
        RECT -4.800 1131.940 2.400 1132.390 ;
        RECT 16.625 1132.375 16.955 1132.390 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 876.420 15.570 876.480 ;
        RECT 610.030 876.420 610.350 876.480 ;
        RECT 15.250 876.280 610.350 876.420 ;
        RECT 15.250 876.220 15.570 876.280 ;
        RECT 610.030 876.220 610.350 876.280 ;
      LAYER via ;
        RECT 15.280 876.220 15.540 876.480 ;
        RECT 610.060 876.220 610.320 876.480 ;
      LAYER met2 ;
        RECT 15.270 881.435 15.550 881.805 ;
        RECT 15.340 876.510 15.480 881.435 ;
        RECT 15.280 876.190 15.540 876.510 ;
        RECT 610.060 876.190 610.320 876.510 ;
        RECT 610.120 855.670 610.260 876.190 ;
        RECT 610.120 855.530 611.640 855.670 ;
        RECT 611.500 749.770 611.640 855.530 ;
        RECT 612.150 749.770 612.430 750.000 ;
        RECT 611.500 749.630 612.430 749.770 ;
        RECT 612.150 746.000 612.430 749.630 ;
      LAYER via2 ;
        RECT 15.270 881.480 15.550 881.760 ;
      LAYER met3 ;
        RECT -4.800 881.770 2.400 882.220 ;
        RECT 15.245 881.770 15.575 881.785 ;
        RECT -4.800 881.470 15.575 881.770 ;
        RECT -4.800 881.020 2.400 881.470 ;
        RECT 15.245 881.455 15.575 881.470 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.550 764.220 615.870 764.280 ;
        RECT 589.420 764.080 615.870 764.220 ;
        RECT 37.790 763.540 38.110 763.600 ;
        RECT 589.420 763.540 589.560 764.080 ;
        RECT 615.550 764.020 615.870 764.080 ;
        RECT 37.790 763.400 589.560 763.540 ;
        RECT 37.790 763.340 38.110 763.400 ;
        RECT 16.630 632.300 16.950 632.360 ;
        RECT 37.790 632.300 38.110 632.360 ;
        RECT 16.630 632.160 38.110 632.300 ;
        RECT 16.630 632.100 16.950 632.160 ;
        RECT 37.790 632.100 38.110 632.160 ;
      LAYER via ;
        RECT 37.820 763.340 38.080 763.600 ;
        RECT 615.580 764.020 615.840 764.280 ;
        RECT 16.660 632.100 16.920 632.360 ;
        RECT 37.820 632.100 38.080 632.360 ;
      LAYER met2 ;
        RECT 615.580 763.990 615.840 764.310 ;
        RECT 37.820 763.310 38.080 763.630 ;
        RECT 37.880 632.390 38.020 763.310 ;
        RECT 615.640 749.770 615.780 763.990 ;
        RECT 616.290 749.770 616.570 750.000 ;
        RECT 615.640 749.630 616.570 749.770 ;
        RECT 616.290 746.000 616.570 749.630 ;
        RECT 16.660 632.070 16.920 632.390 ;
        RECT 37.820 632.070 38.080 632.390 ;
        RECT 16.720 630.885 16.860 632.070 ;
        RECT 16.650 630.515 16.930 630.885 ;
      LAYER via2 ;
        RECT 16.650 630.560 16.930 630.840 ;
      LAYER met3 ;
        RECT -4.800 630.850 2.400 631.300 ;
        RECT 16.625 630.850 16.955 630.865 ;
        RECT -4.800 630.550 16.955 630.850 ;
        RECT -4.800 630.100 2.400 630.550 ;
        RECT 16.625 630.535 16.955 630.550 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 761.840 19.250 761.900 ;
        RECT 619.690 761.840 620.010 761.900 ;
        RECT 18.930 761.700 620.010 761.840 ;
        RECT 18.930 761.640 19.250 761.700 ;
        RECT 619.690 761.640 620.010 761.700 ;
      LAYER via ;
        RECT 18.960 761.640 19.220 761.900 ;
        RECT 619.720 761.640 619.980 761.900 ;
      LAYER met2 ;
        RECT 18.960 761.610 19.220 761.930 ;
        RECT 619.720 761.610 619.980 761.930 ;
        RECT 19.020 379.965 19.160 761.610 ;
        RECT 619.780 749.770 619.920 761.610 ;
        RECT 620.430 749.770 620.710 750.000 ;
        RECT 619.780 749.630 620.710 749.770 ;
        RECT 620.430 746.000 620.710 749.630 ;
        RECT 18.950 379.595 19.230 379.965 ;
      LAYER via2 ;
        RECT 18.950 379.640 19.230 379.920 ;
      LAYER met3 ;
        RECT -4.800 379.930 2.400 380.380 ;
        RECT 18.925 379.930 19.255 379.945 ;
        RECT -4.800 379.630 19.255 379.930 ;
        RECT -4.800 379.180 2.400 379.630 ;
        RECT 18.925 379.615 19.255 379.630 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 755.720 17.870 755.780 ;
        RECT 489.970 755.720 490.290 755.780 ;
        RECT 17.550 755.580 490.290 755.720 ;
        RECT 17.550 755.520 17.870 755.580 ;
        RECT 489.970 755.520 490.290 755.580 ;
      LAYER via ;
        RECT 17.580 755.520 17.840 755.780 ;
        RECT 490.000 755.520 490.260 755.780 ;
      LAYER met2 ;
        RECT 489.990 760.395 490.270 760.765 ;
        RECT 623.850 760.395 624.130 760.765 ;
        RECT 490.060 755.810 490.200 760.395 ;
        RECT 17.580 755.490 17.840 755.810 ;
        RECT 490.000 755.490 490.260 755.810 ;
        RECT 17.640 129.045 17.780 755.490 ;
        RECT 623.920 749.770 624.060 760.395 ;
        RECT 624.570 749.770 624.850 750.000 ;
        RECT 623.920 749.630 624.850 749.770 ;
        RECT 624.570 746.000 624.850 749.630 ;
        RECT 17.570 128.675 17.850 129.045 ;
      LAYER via2 ;
        RECT 489.990 760.440 490.270 760.720 ;
        RECT 623.850 760.440 624.130 760.720 ;
        RECT 17.570 128.720 17.850 129.000 ;
      LAYER met3 ;
        RECT 489.965 760.730 490.295 760.745 ;
        RECT 623.825 760.730 624.155 760.745 ;
        RECT 489.965 760.430 624.155 760.730 ;
        RECT 489.965 760.415 490.295 760.430 ;
        RECT 623.825 760.415 624.155 760.430 ;
        RECT -4.800 129.010 2.400 129.460 ;
        RECT 17.545 129.010 17.875 129.025 ;
        RECT -4.800 128.710 17.875 129.010 ;
        RECT -4.800 128.260 2.400 128.710 ;
        RECT 17.545 128.695 17.875 128.710 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.430 821.340 444.750 821.400 ;
        RECT 2900.830 821.340 2901.150 821.400 ;
        RECT 444.430 821.200 2901.150 821.340 ;
        RECT 444.430 821.140 444.750 821.200 ;
        RECT 2900.830 821.140 2901.150 821.200 ;
      LAYER via ;
        RECT 444.460 821.140 444.720 821.400 ;
        RECT 2900.860 821.140 2901.120 821.400 ;
      LAYER met2 ;
        RECT 444.460 821.110 444.720 821.430 ;
        RECT 2900.860 821.285 2901.120 821.430 ;
        RECT 444.520 749.770 444.660 821.110 ;
        RECT 2900.850 820.915 2901.130 821.285 ;
        RECT 445.170 749.770 445.450 750.000 ;
        RECT 444.520 749.630 445.450 749.770 ;
        RECT 445.170 746.000 445.450 749.630 ;
      LAYER via2 ;
        RECT 2900.850 820.960 2901.130 821.240 ;
      LAYER met3 ;
        RECT 2900.825 821.250 2901.155 821.265 ;
        RECT 2917.600 821.250 2924.800 821.700 ;
        RECT 2900.825 820.950 2924.800 821.250 ;
        RECT 2900.825 820.935 2901.155 820.950 ;
        RECT 2917.600 820.500 2924.800 820.950 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.410 1055.940 450.730 1056.000 ;
        RECT 2900.830 1055.940 2901.150 1056.000 ;
        RECT 450.410 1055.800 2901.150 1055.940 ;
        RECT 450.410 1055.740 450.730 1055.800 ;
        RECT 2900.830 1055.740 2901.150 1055.800 ;
      LAYER via ;
        RECT 450.440 1055.740 450.700 1056.000 ;
        RECT 2900.860 1055.740 2901.120 1056.000 ;
      LAYER met2 ;
        RECT 450.440 1055.710 450.700 1056.030 ;
        RECT 2900.860 1055.885 2901.120 1056.030 ;
        RECT 450.500 751.130 450.640 1055.710 ;
        RECT 2900.850 1055.515 2901.130 1055.885 ;
        RECT 450.500 750.990 450.870 751.130 ;
        RECT 450.730 750.000 450.870 750.990 ;
        RECT 450.690 746.000 450.970 750.000 ;
      LAYER via2 ;
        RECT 2900.850 1055.560 2901.130 1055.840 ;
      LAYER met3 ;
        RECT 2900.825 1055.850 2901.155 1055.865 ;
        RECT 2917.600 1055.850 2924.800 1056.300 ;
        RECT 2900.825 1055.550 2924.800 1055.850 ;
        RECT 2900.825 1055.535 2901.155 1055.550 ;
        RECT 2917.600 1055.100 2924.800 1055.550 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.930 1290.540 456.250 1290.600 ;
        RECT 2904.510 1290.540 2904.830 1290.600 ;
        RECT 455.930 1290.400 2904.830 1290.540 ;
        RECT 455.930 1290.340 456.250 1290.400 ;
        RECT 2904.510 1290.340 2904.830 1290.400 ;
      LAYER via ;
        RECT 455.960 1290.340 456.220 1290.600 ;
        RECT 2904.540 1290.340 2904.800 1290.600 ;
      LAYER met2 ;
        RECT 455.960 1290.310 456.220 1290.630 ;
        RECT 2904.540 1290.485 2904.800 1290.630 ;
        RECT 456.020 751.130 456.160 1290.310 ;
        RECT 2904.530 1290.115 2904.810 1290.485 ;
        RECT 456.020 750.990 456.390 751.130 ;
        RECT 456.250 750.000 456.390 750.990 ;
        RECT 456.210 746.000 456.490 750.000 ;
      LAYER via2 ;
        RECT 2904.530 1290.160 2904.810 1290.440 ;
      LAYER met3 ;
        RECT 2904.505 1290.450 2904.835 1290.465 ;
        RECT 2917.600 1290.450 2924.800 1290.900 ;
        RECT 2904.505 1290.135 2905.050 1290.450 ;
        RECT 2904.750 1289.770 2905.050 1290.135 ;
        RECT 2914.870 1290.150 2924.800 1290.450 ;
        RECT 2914.870 1289.770 2915.170 1290.150 ;
        RECT 2904.750 1289.470 2915.170 1289.770 ;
        RECT 2917.600 1289.700 2924.800 1290.150 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.850 1525.140 457.170 1525.200 ;
        RECT 2900.830 1525.140 2901.150 1525.200 ;
        RECT 456.850 1525.000 2901.150 1525.140 ;
        RECT 456.850 1524.940 457.170 1525.000 ;
        RECT 2900.830 1524.940 2901.150 1525.000 ;
        RECT 456.850 766.600 457.170 766.660 ;
        RECT 460.990 766.600 461.310 766.660 ;
        RECT 456.850 766.460 461.310 766.600 ;
        RECT 456.850 766.400 457.170 766.460 ;
        RECT 460.990 766.400 461.310 766.460 ;
      LAYER via ;
        RECT 456.880 1524.940 457.140 1525.200 ;
        RECT 2900.860 1524.940 2901.120 1525.200 ;
        RECT 456.880 766.400 457.140 766.660 ;
        RECT 461.020 766.400 461.280 766.660 ;
      LAYER met2 ;
        RECT 456.880 1524.910 457.140 1525.230 ;
        RECT 2900.860 1525.085 2901.120 1525.230 ;
        RECT 456.940 766.690 457.080 1524.910 ;
        RECT 2900.850 1524.715 2901.130 1525.085 ;
        RECT 456.880 766.370 457.140 766.690 ;
        RECT 461.020 766.370 461.280 766.690 ;
        RECT 461.080 749.770 461.220 766.370 ;
        RECT 461.730 749.770 462.010 750.000 ;
        RECT 461.080 749.630 462.010 749.770 ;
        RECT 461.730 746.000 462.010 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1524.760 2901.130 1525.040 ;
      LAYER met3 ;
        RECT 2900.825 1525.050 2901.155 1525.065 ;
        RECT 2917.600 1525.050 2924.800 1525.500 ;
        RECT 2900.825 1524.750 2924.800 1525.050 ;
        RECT 2900.825 1524.735 2901.155 1524.750 ;
        RECT 2917.600 1524.300 2924.800 1524.750 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.750 1759.740 464.070 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 463.750 1759.600 2901.150 1759.740 ;
        RECT 463.750 1759.540 464.070 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
        RECT 463.750 796.180 464.070 796.240 ;
        RECT 466.510 796.180 466.830 796.240 ;
        RECT 463.750 796.040 466.830 796.180 ;
        RECT 463.750 795.980 464.070 796.040 ;
        RECT 466.510 795.980 466.830 796.040 ;
      LAYER via ;
        RECT 463.780 1759.540 464.040 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
        RECT 463.780 795.980 464.040 796.240 ;
        RECT 466.540 795.980 466.800 796.240 ;
      LAYER met2 ;
        RECT 463.780 1759.510 464.040 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 463.840 796.270 463.980 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 463.780 795.950 464.040 796.270 ;
        RECT 466.540 795.950 466.800 796.270 ;
        RECT 466.600 749.770 466.740 795.950 ;
        RECT 467.250 749.770 467.530 750.000 ;
        RECT 466.600 749.630 467.530 749.770 ;
        RECT 467.250 746.000 467.530 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.030 1994.340 472.350 1994.400 ;
        RECT 2900.830 1994.340 2901.150 1994.400 ;
        RECT 472.030 1994.200 2901.150 1994.340 ;
        RECT 472.030 1994.140 472.350 1994.200 ;
        RECT 2900.830 1994.140 2901.150 1994.200 ;
      LAYER via ;
        RECT 472.060 1994.140 472.320 1994.400 ;
        RECT 2900.860 1994.140 2901.120 1994.400 ;
      LAYER met2 ;
        RECT 472.060 1994.110 472.320 1994.430 ;
        RECT 2900.860 1994.285 2901.120 1994.430 ;
        RECT 472.120 749.770 472.260 1994.110 ;
        RECT 2900.850 1993.915 2901.130 1994.285 ;
        RECT 472.770 749.770 473.050 750.000 ;
        RECT 472.120 749.630 473.050 749.770 ;
        RECT 472.770 746.000 473.050 749.630 ;
      LAYER via2 ;
        RECT 2900.850 1993.960 2901.130 1994.240 ;
      LAYER met3 ;
        RECT 2900.825 1994.250 2901.155 1994.265 ;
        RECT 2917.600 1994.250 2924.800 1994.700 ;
        RECT 2900.825 1993.950 2924.800 1994.250 ;
        RECT 2900.825 1993.935 2901.155 1993.950 ;
        RECT 2917.600 1993.500 2924.800 1993.950 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.010 2228.940 478.330 2229.000 ;
        RECT 2900.830 2228.940 2901.150 2229.000 ;
        RECT 478.010 2228.800 2901.150 2228.940 ;
        RECT 478.010 2228.740 478.330 2228.800 ;
        RECT 2900.830 2228.740 2901.150 2228.800 ;
      LAYER via ;
        RECT 478.040 2228.740 478.300 2229.000 ;
        RECT 2900.860 2228.740 2901.120 2229.000 ;
      LAYER met2 ;
        RECT 478.040 2228.710 478.300 2229.030 ;
        RECT 2900.860 2228.885 2901.120 2229.030 ;
        RECT 478.100 751.130 478.240 2228.710 ;
        RECT 2900.850 2228.515 2901.130 2228.885 ;
        RECT 478.100 750.990 478.470 751.130 ;
        RECT 478.330 750.000 478.470 750.990 ;
        RECT 478.290 746.000 478.570 750.000 ;
      LAYER via2 ;
        RECT 2900.850 2228.560 2901.130 2228.840 ;
      LAYER met3 ;
        RECT 2900.825 2228.850 2901.155 2228.865 ;
        RECT 2917.600 2228.850 2924.800 2229.300 ;
        RECT 2900.825 2228.550 2924.800 2228.850 ;
        RECT 2900.825 2228.535 2901.155 2228.550 ;
        RECT 2917.600 2228.100 2924.800 2228.550 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 410.390 747.220 410.710 747.280 ;
        RECT 422.810 747.220 423.130 747.280 ;
        RECT 410.390 747.080 423.130 747.220 ;
        RECT 410.390 747.020 410.710 747.080 ;
        RECT 422.810 747.020 423.130 747.080 ;
        RECT 460.760 499.160 461.080 499.420 ;
        RECT 460.070 498.000 460.390 498.060 ;
        RECT 460.850 498.000 460.990 499.160 ;
        RECT 460.070 497.860 460.990 498.000 ;
        RECT 460.070 497.800 460.390 497.860 ;
        RECT 410.390 489.160 410.710 489.220 ;
        RECT 410.390 489.020 460.300 489.160 ;
        RECT 410.390 488.960 410.710 489.020 ;
        RECT 460.160 488.880 460.300 489.020 ;
        RECT 460.070 488.820 460.390 488.880 ;
        RECT 461.910 488.820 462.230 488.880 ;
        RECT 460.070 488.680 462.230 488.820 ;
        RECT 460.070 488.620 460.390 488.680 ;
        RECT 461.910 488.620 462.230 488.680 ;
        RECT 459.150 472.500 459.470 472.560 ;
        RECT 461.910 472.500 462.230 472.560 ;
        RECT 459.150 472.360 462.230 472.500 ;
        RECT 459.150 472.300 459.470 472.360 ;
        RECT 461.910 472.300 462.230 472.360 ;
        RECT 459.150 31.860 459.470 31.920 ;
        RECT 530.910 31.860 531.230 31.920 ;
        RECT 459.150 31.720 531.230 31.860 ;
        RECT 459.150 31.660 459.470 31.720 ;
        RECT 530.910 31.660 531.230 31.720 ;
        RECT 530.910 19.960 531.230 20.020 ;
        RECT 695.130 19.960 695.450 20.020 ;
        RECT 530.910 19.820 695.450 19.960 ;
        RECT 530.910 19.760 531.230 19.820 ;
        RECT 695.130 19.760 695.450 19.820 ;
      LAYER via ;
        RECT 410.420 747.020 410.680 747.280 ;
        RECT 422.840 747.020 423.100 747.280 ;
        RECT 460.790 499.160 461.050 499.420 ;
        RECT 460.100 497.800 460.360 498.060 ;
        RECT 410.420 488.960 410.680 489.220 ;
        RECT 460.100 488.620 460.360 488.880 ;
        RECT 461.940 488.620 462.200 488.880 ;
        RECT 459.180 472.300 459.440 472.560 ;
        RECT 461.940 472.300 462.200 472.560 ;
        RECT 459.180 31.660 459.440 31.920 ;
        RECT 530.940 31.660 531.200 31.920 ;
        RECT 530.940 19.760 531.200 20.020 ;
        RECT 695.160 19.760 695.420 20.020 ;
      LAYER met2 ;
        RECT 410.420 746.990 410.680 747.310 ;
        RECT 422.840 747.050 423.100 747.310 ;
        RECT 424.470 747.050 424.750 750.000 ;
        RECT 422.840 746.990 424.750 747.050 ;
        RECT 410.480 489.250 410.620 746.990 ;
        RECT 422.900 746.910 424.750 746.990 ;
        RECT 424.470 746.000 424.750 746.910 ;
        RECT 460.810 500.000 461.090 504.000 ;
        RECT 460.850 499.450 460.990 500.000 ;
        RECT 460.790 499.130 461.050 499.450 ;
        RECT 460.100 497.770 460.360 498.090 ;
        RECT 410.420 488.930 410.680 489.250 ;
        RECT 460.160 488.910 460.300 497.770 ;
        RECT 460.100 488.590 460.360 488.910 ;
        RECT 461.940 488.590 462.200 488.910 ;
        RECT 462.000 472.590 462.140 488.590 ;
        RECT 459.180 472.270 459.440 472.590 ;
        RECT 461.940 472.270 462.200 472.590 ;
        RECT 459.240 31.950 459.380 472.270 ;
        RECT 459.180 31.630 459.440 31.950 ;
        RECT 530.940 31.630 531.200 31.950 ;
        RECT 531.000 20.050 531.140 31.630 ;
        RECT 530.940 19.730 531.200 20.050 ;
        RECT 695.160 19.730 695.420 20.050 ;
        RECT 695.220 2.400 695.360 19.730 ;
        RECT 695.010 -4.800 695.570 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 492.900 600.690 492.960 ;
        RECT 606.810 492.900 607.130 492.960 ;
        RECT 600.370 492.760 607.130 492.900 ;
        RECT 600.370 492.700 600.690 492.760 ;
        RECT 606.810 492.700 607.130 492.760 ;
        RECT 606.810 487.800 607.130 487.860 ;
        RECT 1003.790 487.800 1004.110 487.860 ;
        RECT 606.810 487.660 1004.110 487.800 ;
        RECT 606.810 487.600 607.130 487.660 ;
        RECT 1003.790 487.600 1004.110 487.660 ;
        RECT 1003.790 440.200 1004.110 440.260 ;
        RECT 2346.070 440.200 2346.390 440.260 ;
        RECT 1003.790 440.060 2346.390 440.200 ;
        RECT 1003.790 440.000 1004.110 440.060 ;
        RECT 2346.070 440.000 2346.390 440.060 ;
      LAYER via ;
        RECT 600.400 492.700 600.660 492.960 ;
        RECT 606.840 492.700 607.100 492.960 ;
        RECT 606.840 487.600 607.100 487.860 ;
        RECT 1003.820 487.600 1004.080 487.860 ;
        RECT 1003.820 440.000 1004.080 440.260 ;
        RECT 2346.100 440.000 2346.360 440.260 ;
      LAYER met2 ;
        RECT 598.810 500.000 599.090 504.000 ;
        RECT 598.850 499.645 598.990 500.000 ;
        RECT 598.780 499.275 599.060 499.645 ;
        RECT 600.390 498.595 600.670 498.965 ;
        RECT 600.460 492.990 600.600 498.595 ;
        RECT 600.400 492.670 600.660 492.990 ;
        RECT 606.840 492.670 607.100 492.990 ;
        RECT 606.900 487.890 607.040 492.670 ;
        RECT 606.840 487.570 607.100 487.890 ;
        RECT 1003.820 487.570 1004.080 487.890 ;
        RECT 1003.880 440.290 1004.020 487.570 ;
        RECT 1003.820 439.970 1004.080 440.290 ;
        RECT 2346.100 439.970 2346.360 440.290 ;
        RECT 2346.160 82.870 2346.300 439.970 ;
        RECT 2346.160 82.730 2351.360 82.870 ;
        RECT 2351.220 2.400 2351.360 82.730 ;
        RECT 2351.010 -4.800 2351.570 2.400 ;
      LAYER via2 ;
        RECT 598.780 499.320 599.060 499.600 ;
        RECT 600.390 498.640 600.670 498.920 ;
      LAYER met3 ;
        RECT 598.755 499.610 599.085 499.625 ;
        RECT 598.755 499.310 600.680 499.610 ;
        RECT 598.755 499.295 599.085 499.310 ;
        RECT 600.380 498.945 600.680 499.310 ;
        RECT 600.365 498.615 600.695 498.945 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.140 499.500 600.460 499.760 ;
        RECT 600.230 498.000 600.370 499.500 ;
        RECT 600.830 498.000 601.150 498.060 ;
        RECT 600.230 497.860 601.150 498.000 ;
        RECT 600.830 497.800 601.150 497.860 ;
        RECT 600.830 470.800 601.150 470.860 ;
        RECT 606.350 470.800 606.670 470.860 ;
        RECT 600.830 470.660 606.670 470.800 ;
        RECT 600.830 470.600 601.150 470.660 ;
        RECT 606.350 470.600 606.670 470.660 ;
        RECT 2367.690 18.260 2368.010 18.320 ;
        RECT 2366.860 18.120 2368.010 18.260 ;
        RECT 606.350 17.920 606.670 17.980 ;
        RECT 2366.860 17.920 2367.000 18.120 ;
        RECT 2367.690 18.060 2368.010 18.120 ;
        RECT 606.350 17.780 2367.000 17.920 ;
        RECT 606.350 17.720 606.670 17.780 ;
      LAYER via ;
        RECT 600.170 499.500 600.430 499.760 ;
        RECT 600.860 497.800 601.120 498.060 ;
        RECT 600.860 470.600 601.120 470.860 ;
        RECT 606.380 470.600 606.640 470.860 ;
        RECT 606.380 17.720 606.640 17.980 ;
        RECT 2367.720 18.060 2367.980 18.320 ;
      LAYER met2 ;
        RECT 600.190 500.000 600.470 504.000 ;
        RECT 600.230 499.790 600.370 500.000 ;
        RECT 600.170 499.470 600.430 499.790 ;
        RECT 600.860 497.770 601.120 498.090 ;
        RECT 600.920 470.890 601.060 497.770 ;
        RECT 600.860 470.570 601.120 470.890 ;
        RECT 606.380 470.570 606.640 470.890 ;
        RECT 606.440 18.010 606.580 470.570 ;
        RECT 2367.720 18.030 2367.980 18.350 ;
        RECT 606.380 17.690 606.640 18.010 ;
        RECT 2367.780 2.400 2367.920 18.030 ;
        RECT 2367.570 -4.800 2368.130 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 483.720 602.070 483.780 ;
        RECT 639.930 483.720 640.250 483.780 ;
        RECT 601.750 483.580 640.250 483.720 ;
        RECT 601.750 483.520 602.070 483.580 ;
        RECT 639.930 483.520 640.250 483.580 ;
        RECT 2384.250 18.600 2384.570 18.660 ;
        RECT 2352.830 18.460 2384.570 18.600 ;
        RECT 639.930 18.260 640.250 18.320 ;
        RECT 2352.830 18.260 2352.970 18.460 ;
        RECT 2384.250 18.400 2384.570 18.460 ;
        RECT 639.930 18.120 2352.970 18.260 ;
        RECT 639.930 18.060 640.250 18.120 ;
      LAYER via ;
        RECT 601.780 483.520 602.040 483.780 ;
        RECT 639.960 483.520 640.220 483.780 ;
        RECT 639.960 18.060 640.220 18.320 ;
        RECT 2384.280 18.400 2384.540 18.660 ;
      LAYER met2 ;
        RECT 601.570 500.000 601.850 504.000 ;
        RECT 601.610 499.020 601.750 500.000 ;
        RECT 601.610 498.880 601.980 499.020 ;
        RECT 601.840 498.680 601.980 498.880 ;
        RECT 601.840 498.540 602.210 498.680 ;
        RECT 602.070 498.170 602.210 498.540 ;
        RECT 601.840 498.030 602.210 498.170 ;
        RECT 601.840 483.810 601.980 498.030 ;
        RECT 601.780 483.490 602.040 483.810 ;
        RECT 639.960 483.490 640.220 483.810 ;
        RECT 640.020 18.350 640.160 483.490 ;
        RECT 2384.280 18.370 2384.540 18.690 ;
        RECT 639.960 18.030 640.220 18.350 ;
        RECT 2384.340 2.400 2384.480 18.370 ;
        RECT 2384.130 -4.800 2384.690 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 602.900 499.500 603.220 499.760 ;
        RECT 602.990 499.020 603.130 499.500 ;
        RECT 602.990 498.880 603.360 499.020 ;
        RECT 603.220 498.740 603.360 498.880 ;
        RECT 603.130 498.480 603.450 498.740 ;
        RECT 603.590 176.360 603.910 176.420 ;
        RECT 2394.370 176.360 2394.690 176.420 ;
        RECT 603.590 176.220 2394.690 176.360 ;
        RECT 603.590 176.160 603.910 176.220 ;
        RECT 2394.370 176.160 2394.690 176.220 ;
        RECT 2394.370 5.680 2394.690 5.740 ;
        RECT 2400.810 5.680 2401.130 5.740 ;
        RECT 2394.370 5.540 2401.130 5.680 ;
        RECT 2394.370 5.480 2394.690 5.540 ;
        RECT 2400.810 5.480 2401.130 5.540 ;
      LAYER via ;
        RECT 602.930 499.500 603.190 499.760 ;
        RECT 603.160 498.480 603.420 498.740 ;
        RECT 603.620 176.160 603.880 176.420 ;
        RECT 2394.400 176.160 2394.660 176.420 ;
        RECT 2394.400 5.480 2394.660 5.740 ;
        RECT 2400.840 5.480 2401.100 5.740 ;
      LAYER met2 ;
        RECT 602.950 500.000 603.230 504.000 ;
        RECT 602.990 499.790 603.130 500.000 ;
        RECT 602.930 499.470 603.190 499.790 ;
        RECT 603.160 498.450 603.420 498.770 ;
        RECT 603.220 485.250 603.360 498.450 ;
        RECT 603.220 485.110 603.820 485.250 ;
        RECT 603.680 176.450 603.820 485.110 ;
        RECT 603.620 176.130 603.880 176.450 ;
        RECT 2394.400 176.130 2394.660 176.450 ;
        RECT 2394.460 5.770 2394.600 176.130 ;
        RECT 2394.400 5.450 2394.660 5.770 ;
        RECT 2400.840 5.450 2401.100 5.770 ;
        RECT 2400.900 2.400 2401.040 5.450 ;
        RECT 2400.690 -4.800 2401.250 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.050 484.740 604.370 484.800 ;
        RECT 604.970 484.740 605.290 484.800 ;
        RECT 604.050 484.600 605.290 484.740 ;
        RECT 604.050 484.540 604.370 484.600 ;
        RECT 604.970 484.540 605.290 484.600 ;
        RECT 604.050 197.440 604.370 197.500 ;
        RECT 2415.070 197.440 2415.390 197.500 ;
        RECT 604.050 197.300 2415.390 197.440 ;
        RECT 604.050 197.240 604.370 197.300 ;
        RECT 2415.070 197.240 2415.390 197.300 ;
      LAYER via ;
        RECT 604.080 484.540 604.340 484.800 ;
        RECT 605.000 484.540 605.260 484.800 ;
        RECT 604.080 197.240 604.340 197.500 ;
        RECT 2415.100 197.240 2415.360 197.500 ;
      LAYER met2 ;
        RECT 604.330 500.000 604.610 504.000 ;
        RECT 604.370 498.850 604.510 500.000 ;
        RECT 604.370 498.710 604.740 498.850 ;
        RECT 604.600 485.760 604.740 498.710 ;
        RECT 604.600 485.620 605.200 485.760 ;
        RECT 605.060 484.830 605.200 485.620 ;
        RECT 604.080 484.510 604.340 484.830 ;
        RECT 605.000 484.510 605.260 484.830 ;
        RECT 604.140 197.530 604.280 484.510 ;
        RECT 604.080 197.210 604.340 197.530 ;
        RECT 2415.100 197.210 2415.360 197.530 ;
        RECT 2415.160 82.870 2415.300 197.210 ;
        RECT 2415.160 82.730 2417.600 82.870 ;
        RECT 2417.460 2.400 2417.600 82.730 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.710 500.000 605.990 504.000 ;
        RECT 605.750 499.020 605.890 500.000 ;
        RECT 605.520 498.880 605.890 499.020 ;
        RECT 605.520 498.850 605.660 498.880 ;
        RECT 605.290 498.710 605.660 498.850 ;
        RECT 605.290 498.170 605.430 498.710 ;
        RECT 605.290 498.030 605.660 498.170 ;
        RECT 605.520 486.045 605.660 498.030 ;
        RECT 605.450 485.675 605.730 486.045 ;
        RECT 2428.890 452.355 2429.170 452.725 ;
        RECT 2428.960 82.870 2429.100 452.355 ;
        RECT 2428.960 82.730 2434.160 82.870 ;
        RECT 2434.020 2.400 2434.160 82.730 ;
        RECT 2433.810 -4.800 2434.370 2.400 ;
      LAYER via2 ;
        RECT 605.450 485.720 605.730 486.000 ;
        RECT 2428.890 452.400 2429.170 452.680 ;
      LAYER met3 ;
        RECT 602.870 486.010 603.250 486.020 ;
        RECT 605.425 486.010 605.755 486.025 ;
        RECT 602.870 485.710 605.755 486.010 ;
        RECT 602.870 485.700 603.250 485.710 ;
        RECT 605.425 485.695 605.755 485.710 ;
        RECT 602.870 452.690 603.250 452.700 ;
        RECT 2428.865 452.690 2429.195 452.705 ;
        RECT 602.870 452.390 2429.195 452.690 ;
        RECT 602.870 452.380 603.250 452.390 ;
        RECT 2428.865 452.375 2429.195 452.390 ;
      LAYER via3 ;
        RECT 602.900 485.700 603.220 486.020 ;
        RECT 602.900 452.380 603.220 452.700 ;
      LAYER met4 ;
        RECT 602.895 485.695 603.225 486.025 ;
        RECT 602.910 452.705 603.210 485.695 ;
        RECT 602.895 452.375 603.225 452.705 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.040 499.700 607.360 499.760 ;
        RECT 607.040 499.560 610.720 499.700 ;
        RECT 607.040 499.500 607.360 499.560 ;
        RECT 610.580 497.660 610.720 499.560 ;
        RECT 610.580 497.520 613.020 497.660 ;
        RECT 612.880 497.320 613.020 497.520 ;
        RECT 613.710 497.320 614.030 497.380 ;
        RECT 612.880 497.180 614.030 497.320 ;
        RECT 613.710 497.120 614.030 497.180 ;
        RECT 613.710 487.120 614.030 487.180 ;
        RECT 1390.190 487.120 1390.510 487.180 ;
        RECT 613.710 486.980 1390.510 487.120 ;
        RECT 613.710 486.920 614.030 486.980 ;
        RECT 1390.190 486.920 1390.510 486.980 ;
        RECT 1390.190 19.960 1390.510 20.020 ;
        RECT 1390.190 19.820 1435.270 19.960 ;
        RECT 1390.190 19.760 1390.510 19.820 ;
        RECT 1435.130 19.620 1435.270 19.820 ;
        RECT 2450.490 19.620 2450.810 19.680 ;
        RECT 1435.130 19.480 2450.810 19.620 ;
        RECT 2450.490 19.420 2450.810 19.480 ;
      LAYER via ;
        RECT 607.070 499.500 607.330 499.760 ;
        RECT 613.740 497.120 614.000 497.380 ;
        RECT 613.740 486.920 614.000 487.180 ;
        RECT 1390.220 486.920 1390.480 487.180 ;
        RECT 1390.220 19.760 1390.480 20.020 ;
        RECT 2450.520 19.420 2450.780 19.680 ;
      LAYER met2 ;
        RECT 607.090 500.000 607.370 504.000 ;
        RECT 607.130 499.790 607.270 500.000 ;
        RECT 607.070 499.470 607.330 499.790 ;
        RECT 613.740 497.090 614.000 497.410 ;
        RECT 613.800 487.210 613.940 497.090 ;
        RECT 613.740 486.890 614.000 487.210 ;
        RECT 1390.220 486.890 1390.480 487.210 ;
        RECT 1390.280 20.050 1390.420 486.890 ;
        RECT 1390.220 19.730 1390.480 20.050 ;
        RECT 2450.520 19.390 2450.780 19.710 ;
        RECT 2450.580 2.400 2450.720 19.390 ;
        RECT 2450.370 -4.800 2450.930 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 474.880 608.510 474.940 ;
        RECT 612.790 474.880 613.110 474.940 ;
        RECT 608.190 474.740 613.110 474.880 ;
        RECT 608.190 474.680 608.510 474.740 ;
        RECT 612.790 474.680 613.110 474.740 ;
        RECT 2467.050 17.920 2467.370 17.980 ;
        RECT 2449.430 17.780 2467.370 17.920 ;
        RECT 612.790 17.580 613.110 17.640 ;
        RECT 2449.430 17.580 2449.570 17.780 ;
        RECT 2467.050 17.720 2467.370 17.780 ;
        RECT 612.790 17.440 2449.570 17.580 ;
        RECT 612.790 17.380 613.110 17.440 ;
      LAYER via ;
        RECT 608.220 474.680 608.480 474.940 ;
        RECT 612.820 474.680 613.080 474.940 ;
        RECT 612.820 17.380 613.080 17.640 ;
        RECT 2467.080 17.720 2467.340 17.980 ;
      LAYER met2 ;
        RECT 608.470 500.000 608.750 504.000 ;
        RECT 608.510 499.475 608.650 500.000 ;
        RECT 608.440 499.105 608.720 499.475 ;
        RECT 608.210 497.915 608.490 498.285 ;
        RECT 608.280 474.970 608.420 497.915 ;
        RECT 608.220 474.650 608.480 474.970 ;
        RECT 612.820 474.650 613.080 474.970 ;
        RECT 612.880 17.670 613.020 474.650 ;
        RECT 2467.080 17.690 2467.340 18.010 ;
        RECT 612.820 17.350 613.080 17.670 ;
        RECT 2467.140 2.400 2467.280 17.690 ;
        RECT 2466.930 -4.800 2467.490 2.400 ;
      LAYER via2 ;
        RECT 608.440 499.150 608.720 499.430 ;
        RECT 608.210 497.960 608.490 498.240 ;
      LAYER met3 ;
        RECT 608.415 499.125 608.745 499.455 ;
        RECT 608.430 498.265 608.730 499.125 ;
        RECT 608.185 497.950 608.730 498.265 ;
        RECT 608.185 497.935 608.515 497.950 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 476.920 608.050 476.980 ;
        RECT 609.570 476.920 609.890 476.980 ;
        RECT 607.730 476.780 609.890 476.920 ;
        RECT 607.730 476.720 608.050 476.780 ;
        RECT 609.570 476.720 609.890 476.780 ;
        RECT 607.730 17.240 608.050 17.300 ;
        RECT 2483.610 17.240 2483.930 17.300 ;
        RECT 607.730 17.100 2483.930 17.240 ;
        RECT 607.730 17.040 608.050 17.100 ;
        RECT 2483.610 17.040 2483.930 17.100 ;
      LAYER via ;
        RECT 607.760 476.720 608.020 476.980 ;
        RECT 609.600 476.720 609.860 476.980 ;
        RECT 607.760 17.040 608.020 17.300 ;
        RECT 2483.640 17.040 2483.900 17.300 ;
      LAYER met2 ;
        RECT 609.850 500.000 610.130 504.000 ;
        RECT 609.890 498.850 610.030 500.000 ;
        RECT 609.660 498.710 610.030 498.850 ;
        RECT 609.660 477.010 609.800 498.710 ;
        RECT 607.760 476.690 608.020 477.010 ;
        RECT 609.600 476.690 609.860 477.010 ;
        RECT 607.820 17.330 607.960 476.690 ;
        RECT 607.760 17.010 608.020 17.330 ;
        RECT 2483.640 17.010 2483.900 17.330 ;
        RECT 2483.700 2.400 2483.840 17.010 ;
        RECT 2483.490 -4.800 2484.050 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.180 499.500 611.500 499.760 ;
        RECT 611.270 498.340 611.410 499.500 ;
        RECT 611.870 498.340 612.190 498.400 ;
        RECT 611.270 498.200 612.190 498.340 ;
        RECT 611.870 498.140 612.190 498.200 ;
        RECT 608.190 471.480 608.510 471.540 ;
        RECT 611.870 471.480 612.190 471.540 ;
        RECT 608.190 471.340 612.190 471.480 ;
        RECT 608.190 471.280 608.510 471.340 ;
        RECT 611.870 471.280 612.190 471.340 ;
        RECT 608.190 25.400 608.510 25.460 ;
        RECT 2500.170 25.400 2500.490 25.460 ;
        RECT 608.190 25.260 2500.490 25.400 ;
        RECT 608.190 25.200 608.510 25.260 ;
        RECT 2500.170 25.200 2500.490 25.260 ;
      LAYER via ;
        RECT 611.210 499.500 611.470 499.760 ;
        RECT 611.900 498.140 612.160 498.400 ;
        RECT 608.220 471.280 608.480 471.540 ;
        RECT 611.900 471.280 612.160 471.540 ;
        RECT 608.220 25.200 608.480 25.460 ;
        RECT 2500.200 25.200 2500.460 25.460 ;
      LAYER met2 ;
        RECT 611.230 500.000 611.510 504.000 ;
        RECT 611.270 499.790 611.410 500.000 ;
        RECT 611.210 499.470 611.470 499.790 ;
        RECT 611.900 498.110 612.160 498.430 ;
        RECT 611.960 471.570 612.100 498.110 ;
        RECT 608.220 471.250 608.480 471.570 ;
        RECT 611.900 471.250 612.160 471.570 ;
        RECT 608.280 25.490 608.420 471.250 ;
        RECT 608.220 25.170 608.480 25.490 ;
        RECT 2500.200 25.170 2500.460 25.490 ;
        RECT 2500.260 2.400 2500.400 25.170 ;
        RECT 2500.050 -4.800 2500.610 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 409.470 762.860 409.790 762.920 ;
        RECT 478.930 762.860 479.250 762.920 ;
        RECT 409.470 762.720 479.250 762.860 ;
        RECT 409.470 762.660 409.790 762.720 ;
        RECT 478.930 762.660 479.250 762.720 ;
        RECT 409.010 501.400 409.330 501.460 ;
        RECT 409.010 501.260 464.210 501.400 ;
        RECT 409.010 501.200 409.330 501.260 ;
        RECT 464.070 501.060 464.210 501.260 ;
        RECT 464.070 500.920 474.790 501.060 ;
        RECT 474.650 499.760 474.790 500.920 ;
        RECT 474.560 499.500 474.880 499.760 ;
        RECT 474.650 499.020 474.790 499.500 ;
        RECT 474.650 498.880 475.020 499.020 ;
        RECT 474.880 498.400 475.020 498.880 ;
        RECT 474.790 498.140 475.110 498.400 ;
        RECT 474.790 486.100 475.110 486.160 ;
        RECT 474.790 485.960 496.870 486.100 ;
        RECT 474.790 485.900 475.110 485.960 ;
        RECT 496.730 483.380 496.870 485.960 ;
        RECT 606.810 483.380 607.130 483.440 ;
        RECT 496.730 483.240 607.130 483.380 ;
        RECT 606.810 483.180 607.130 483.240 ;
        RECT 606.810 461.620 607.130 461.680 ;
        RECT 855.670 461.620 855.990 461.680 ;
        RECT 606.810 461.480 855.990 461.620 ;
        RECT 606.810 461.420 607.130 461.480 ;
        RECT 855.670 461.420 855.990 461.480 ;
      LAYER via ;
        RECT 409.500 762.660 409.760 762.920 ;
        RECT 478.960 762.660 479.220 762.920 ;
        RECT 409.040 501.200 409.300 501.460 ;
        RECT 474.590 499.500 474.850 499.760 ;
        RECT 474.820 498.140 475.080 498.400 ;
        RECT 474.820 485.900 475.080 486.160 ;
        RECT 606.840 483.180 607.100 483.440 ;
        RECT 606.840 461.420 607.100 461.680 ;
        RECT 855.700 461.420 855.960 461.680 ;
      LAYER met2 ;
        RECT 409.500 762.630 409.760 762.950 ;
        RECT 478.960 762.630 479.220 762.950 ;
        RECT 409.560 521.290 409.700 762.630 ;
        RECT 479.020 749.770 479.160 762.630 ;
        RECT 479.670 749.770 479.950 750.000 ;
        RECT 479.020 749.630 479.950 749.770 ;
        RECT 479.670 746.000 479.950 749.630 ;
        RECT 409.100 521.150 409.700 521.290 ;
        RECT 409.100 501.490 409.240 521.150 ;
        RECT 409.040 501.170 409.300 501.490 ;
        RECT 474.610 500.000 474.890 504.000 ;
        RECT 474.650 499.790 474.790 500.000 ;
        RECT 474.590 499.470 474.850 499.790 ;
        RECT 474.820 498.110 475.080 498.430 ;
        RECT 474.880 486.190 475.020 498.110 ;
        RECT 474.820 485.870 475.080 486.190 ;
        RECT 606.840 483.150 607.100 483.470 ;
        RECT 606.900 461.710 607.040 483.150 ;
        RECT 606.840 461.390 607.100 461.710 ;
        RECT 855.700 461.390 855.960 461.710 ;
        RECT 855.760 82.870 855.900 461.390 ;
        RECT 855.760 82.730 860.960 82.870 ;
        RECT 860.820 2.400 860.960 82.730 ;
        RECT 860.610 -4.800 861.170 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.610 500.000 612.890 504.000 ;
        RECT 612.650 499.645 612.790 500.000 ;
        RECT 612.580 499.275 612.860 499.645 ;
        RECT 2511.690 451.675 2511.970 452.045 ;
        RECT 2511.760 82.870 2511.900 451.675 ;
        RECT 2511.760 82.730 2516.960 82.870 ;
        RECT 2516.820 2.400 2516.960 82.730 ;
        RECT 2516.610 -4.800 2517.170 2.400 ;
      LAYER via2 ;
        RECT 612.580 499.320 612.860 499.600 ;
        RECT 2511.690 451.720 2511.970 452.000 ;
      LAYER met3 ;
        RECT 612.555 499.610 612.885 499.625 ;
        RECT 612.555 499.295 613.100 499.610 ;
        RECT 612.800 498.940 613.100 499.295 ;
        RECT 612.800 498.630 613.370 498.940 ;
        RECT 612.990 498.620 613.370 498.630 ;
        RECT 612.990 452.010 613.370 452.020 ;
        RECT 2511.665 452.010 2511.995 452.025 ;
        RECT 612.990 451.710 2511.995 452.010 ;
        RECT 612.990 451.700 613.370 451.710 ;
        RECT 2511.665 451.695 2511.995 451.710 ;
      LAYER via3 ;
        RECT 613.020 498.620 613.340 498.940 ;
        RECT 613.020 451.700 613.340 452.020 ;
      LAYER met4 ;
        RECT 613.015 498.615 613.345 498.945 ;
        RECT 613.030 452.025 613.330 498.615 ;
        RECT 613.015 451.695 613.345 452.025 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.940 499.840 614.260 500.100 ;
        RECT 614.030 497.660 614.170 499.840 ;
        RECT 617.850 497.660 618.170 497.720 ;
        RECT 614.030 497.520 618.170 497.660 ;
        RECT 617.850 497.460 618.170 497.520 ;
        RECT 617.850 483.380 618.170 483.440 ;
        RECT 625.670 483.380 625.990 483.440 ;
        RECT 617.850 483.240 625.990 483.380 ;
        RECT 617.850 483.180 618.170 483.240 ;
        RECT 625.670 483.180 625.990 483.240 ;
        RECT 625.670 458.900 625.990 458.960 ;
        RECT 2532.370 458.900 2532.690 458.960 ;
        RECT 625.670 458.760 2532.690 458.900 ;
        RECT 625.670 458.700 625.990 458.760 ;
        RECT 2532.370 458.700 2532.690 458.760 ;
      LAYER via ;
        RECT 613.970 499.840 614.230 500.100 ;
        RECT 617.880 497.460 618.140 497.720 ;
        RECT 617.880 483.180 618.140 483.440 ;
        RECT 625.700 483.180 625.960 483.440 ;
        RECT 625.700 458.700 625.960 458.960 ;
        RECT 2532.400 458.700 2532.660 458.960 ;
      LAYER met2 ;
        RECT 613.990 500.130 614.270 504.000 ;
        RECT 613.970 500.000 614.270 500.130 ;
        RECT 613.970 499.810 614.230 500.000 ;
        RECT 617.880 497.430 618.140 497.750 ;
        RECT 617.940 483.470 618.080 497.430 ;
        RECT 617.880 483.150 618.140 483.470 ;
        RECT 625.700 483.150 625.960 483.470 ;
        RECT 625.760 458.990 625.900 483.150 ;
        RECT 625.700 458.670 625.960 458.990 ;
        RECT 2532.400 458.670 2532.660 458.990 ;
        RECT 2532.460 17.410 2532.600 458.670 ;
        RECT 2532.460 17.270 2533.520 17.410 ;
        RECT 2533.380 2.400 2533.520 17.270 ;
        RECT 2533.170 -4.800 2533.730 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.320 499.160 615.640 499.420 ;
        RECT 614.630 498.340 614.950 498.400 ;
        RECT 615.410 498.340 615.550 499.160 ;
        RECT 614.630 498.200 615.550 498.340 ;
        RECT 614.630 498.140 614.950 498.200 ;
        RECT 614.170 25.060 614.490 25.120 ;
        RECT 2549.850 25.060 2550.170 25.120 ;
        RECT 614.170 24.920 2550.170 25.060 ;
        RECT 614.170 24.860 614.490 24.920 ;
        RECT 2549.850 24.860 2550.170 24.920 ;
      LAYER via ;
        RECT 615.350 499.160 615.610 499.420 ;
        RECT 614.660 498.140 614.920 498.400 ;
        RECT 614.200 24.860 614.460 25.120 ;
        RECT 2549.880 24.860 2550.140 25.120 ;
      LAYER met2 ;
        RECT 615.370 500.000 615.650 504.000 ;
        RECT 615.410 499.450 615.550 500.000 ;
        RECT 615.350 499.130 615.610 499.450 ;
        RECT 614.660 498.110 614.920 498.430 ;
        RECT 614.720 473.010 614.860 498.110 ;
        RECT 614.260 472.870 614.860 473.010 ;
        RECT 614.260 25.150 614.400 472.870 ;
        RECT 614.200 24.830 614.460 25.150 ;
        RECT 2549.880 24.830 2550.140 25.150 ;
        RECT 2549.940 2.400 2550.080 24.830 ;
        RECT 2549.730 -4.800 2550.290 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.850 439.180 618.170 439.240 ;
        RECT 2559.970 439.180 2560.290 439.240 ;
        RECT 617.850 439.040 2560.290 439.180 ;
        RECT 617.850 438.980 618.170 439.040 ;
        RECT 2559.970 438.980 2560.290 439.040 ;
        RECT 2559.970 17.580 2560.290 17.640 ;
        RECT 2566.410 17.580 2566.730 17.640 ;
        RECT 2559.970 17.440 2566.730 17.580 ;
        RECT 2559.970 17.380 2560.290 17.440 ;
        RECT 2566.410 17.380 2566.730 17.440 ;
      LAYER via ;
        RECT 617.880 438.980 618.140 439.240 ;
        RECT 2560.000 438.980 2560.260 439.240 ;
        RECT 2560.000 17.380 2560.260 17.640 ;
        RECT 2566.440 17.380 2566.700 17.640 ;
      LAYER met2 ;
        RECT 616.750 500.000 617.030 504.000 ;
        RECT 616.790 499.020 616.930 500.000 ;
        RECT 616.790 498.880 617.620 499.020 ;
        RECT 617.480 475.730 617.620 498.880 ;
        RECT 617.480 475.590 618.080 475.730 ;
        RECT 617.940 439.270 618.080 475.590 ;
        RECT 617.880 438.950 618.140 439.270 ;
        RECT 2560.000 438.950 2560.260 439.270 ;
        RECT 2560.060 17.670 2560.200 438.950 ;
        RECT 2560.000 17.350 2560.260 17.670 ;
        RECT 2566.440 17.350 2566.700 17.670 ;
        RECT 2566.500 2.400 2566.640 17.350 ;
        RECT 2566.290 -4.800 2566.850 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.310 438.840 618.630 438.900 ;
        RECT 2580.670 438.840 2580.990 438.900 ;
        RECT 618.310 438.700 2580.990 438.840 ;
        RECT 618.310 438.640 618.630 438.700 ;
        RECT 2580.670 438.640 2580.990 438.700 ;
      LAYER via ;
        RECT 618.340 438.640 618.600 438.900 ;
        RECT 2580.700 438.640 2580.960 438.900 ;
      LAYER met2 ;
        RECT 618.130 500.000 618.410 504.000 ;
        RECT 618.170 498.850 618.310 500.000 ;
        RECT 618.170 498.710 618.540 498.850 ;
        RECT 618.400 438.930 618.540 498.710 ;
        RECT 618.340 438.610 618.600 438.930 ;
        RECT 2580.700 438.610 2580.960 438.930 ;
        RECT 2580.760 82.870 2580.900 438.610 ;
        RECT 2580.760 82.730 2583.200 82.870 ;
        RECT 2583.060 2.400 2583.200 82.730 ;
        RECT 2582.850 -4.800 2583.410 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.510 500.000 619.790 504.000 ;
        RECT 619.550 499.645 619.690 500.000 ;
        RECT 619.480 499.275 619.760 499.645 ;
        RECT 2599.550 23.955 2599.830 24.325 ;
        RECT 2599.620 2.400 2599.760 23.955 ;
        RECT 2599.410 -4.800 2599.970 2.400 ;
      LAYER via2 ;
        RECT 619.480 499.320 619.760 499.600 ;
        RECT 2599.550 24.000 2599.830 24.280 ;
      LAYER met3 ;
        RECT 619.455 499.610 619.785 499.625 ;
        RECT 620.350 499.610 620.730 499.620 ;
        RECT 619.455 499.310 620.730 499.610 ;
        RECT 619.455 499.295 619.785 499.310 ;
        RECT 620.350 499.300 620.730 499.310 ;
        RECT 620.350 24.290 620.730 24.300 ;
        RECT 2599.525 24.290 2599.855 24.305 ;
        RECT 620.350 23.990 2599.855 24.290 ;
        RECT 620.350 23.980 620.730 23.990 ;
        RECT 2599.525 23.975 2599.855 23.990 ;
      LAYER via3 ;
        RECT 620.380 499.300 620.700 499.620 ;
        RECT 620.380 23.980 620.700 24.300 ;
      LAYER met4 ;
        RECT 620.375 499.295 620.705 499.625 ;
        RECT 620.390 24.305 620.690 499.295 ;
        RECT 620.375 23.975 620.705 24.305 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 620.840 499.160 621.160 499.420 ;
        RECT 620.930 498.340 621.070 499.160 ;
        RECT 622.450 498.340 622.770 498.400 ;
        RECT 620.930 498.200 622.770 498.340 ;
        RECT 622.450 498.140 622.770 498.200 ;
        RECT 622.450 486.440 622.770 486.500 ;
        RECT 2231.990 486.440 2232.310 486.500 ;
        RECT 622.450 486.300 2232.310 486.440 ;
        RECT 622.450 486.240 622.770 486.300 ;
        RECT 2231.990 486.240 2232.310 486.300 ;
        RECT 2231.990 19.280 2232.310 19.340 ;
        RECT 2231.990 19.140 2256.370 19.280 ;
        RECT 2231.990 19.080 2232.310 19.140 ;
        RECT 2256.230 18.940 2256.370 19.140 ;
        RECT 2616.090 18.940 2616.410 19.000 ;
        RECT 2256.230 18.800 2616.410 18.940 ;
        RECT 2616.090 18.740 2616.410 18.800 ;
      LAYER via ;
        RECT 620.870 499.160 621.130 499.420 ;
        RECT 622.480 498.140 622.740 498.400 ;
        RECT 622.480 486.240 622.740 486.500 ;
        RECT 2232.020 486.240 2232.280 486.500 ;
        RECT 2232.020 19.080 2232.280 19.340 ;
        RECT 2616.120 18.740 2616.380 19.000 ;
      LAYER met2 ;
        RECT 620.890 500.000 621.170 504.000 ;
        RECT 620.930 499.450 621.070 500.000 ;
        RECT 620.870 499.130 621.130 499.450 ;
        RECT 622.480 498.110 622.740 498.430 ;
        RECT 622.540 486.530 622.680 498.110 ;
        RECT 622.480 486.210 622.740 486.530 ;
        RECT 2232.020 486.210 2232.280 486.530 ;
        RECT 2232.080 19.370 2232.220 486.210 ;
        RECT 2232.020 19.050 2232.280 19.370 ;
        RECT 2616.120 18.710 2616.380 19.030 ;
        RECT 2616.180 2.400 2616.320 18.710 ;
        RECT 2615.970 -4.800 2616.530 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.530 498.680 621.850 498.740 ;
        RECT 621.990 498.680 622.310 498.740 ;
        RECT 621.530 498.540 622.310 498.680 ;
        RECT 621.530 498.480 621.850 498.540 ;
        RECT 621.990 498.480 622.310 498.540 ;
        RECT 621.530 24.720 621.850 24.780 ;
        RECT 2632.650 24.720 2632.970 24.780 ;
        RECT 621.530 24.580 2632.970 24.720 ;
        RECT 621.530 24.520 621.850 24.580 ;
        RECT 2632.650 24.520 2632.970 24.580 ;
      LAYER via ;
        RECT 621.560 498.480 621.820 498.740 ;
        RECT 622.020 498.480 622.280 498.740 ;
        RECT 621.560 24.520 621.820 24.780 ;
        RECT 2632.680 24.520 2632.940 24.780 ;
      LAYER met2 ;
        RECT 622.270 500.000 622.550 504.000 ;
        RECT 622.310 498.850 622.450 500.000 ;
        RECT 622.080 498.770 622.450 498.850 ;
        RECT 621.560 498.450 621.820 498.770 ;
        RECT 622.020 498.710 622.450 498.770 ;
        RECT 622.020 498.450 622.280 498.710 ;
        RECT 621.620 24.810 621.760 498.450 ;
        RECT 621.560 24.490 621.820 24.810 ;
        RECT 2632.680 24.490 2632.940 24.810 ;
        RECT 2632.740 2.400 2632.880 24.490 ;
        RECT 2632.530 -4.800 2633.090 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 623.600 500.040 623.920 500.100 ;
        RECT 623.600 499.840 624.060 500.040 ;
        RECT 621.070 497.660 621.390 497.720 ;
        RECT 623.920 497.660 624.060 499.840 ;
        RECT 621.070 497.520 624.060 497.660 ;
        RECT 621.070 497.460 621.390 497.520 ;
        RECT 621.070 24.380 621.390 24.440 ;
        RECT 2583.890 24.380 2584.210 24.440 ;
        RECT 621.070 24.240 2584.210 24.380 ;
        RECT 621.070 24.180 621.390 24.240 ;
        RECT 2583.890 24.180 2584.210 24.240 ;
        RECT 2583.890 23.700 2584.210 23.760 ;
        RECT 2649.210 23.700 2649.530 23.760 ;
        RECT 2583.890 23.560 2649.530 23.700 ;
        RECT 2583.890 23.500 2584.210 23.560 ;
        RECT 2649.210 23.500 2649.530 23.560 ;
      LAYER via ;
        RECT 623.630 499.840 623.890 500.100 ;
        RECT 621.100 497.460 621.360 497.720 ;
        RECT 621.100 24.180 621.360 24.440 ;
        RECT 2583.920 24.180 2584.180 24.440 ;
        RECT 2583.920 23.500 2584.180 23.760 ;
        RECT 2649.240 23.500 2649.500 23.760 ;
      LAYER met2 ;
        RECT 623.650 500.130 623.930 504.000 ;
        RECT 623.630 500.000 623.930 500.130 ;
        RECT 623.630 499.810 623.890 500.000 ;
        RECT 621.100 497.430 621.360 497.750 ;
        RECT 621.160 24.470 621.300 497.430 ;
        RECT 621.100 24.150 621.360 24.470 ;
        RECT 2583.920 24.150 2584.180 24.470 ;
        RECT 2583.980 23.790 2584.120 24.150 ;
        RECT 2583.920 23.470 2584.180 23.790 ;
        RECT 2649.240 23.470 2649.500 23.790 ;
        RECT 2649.300 2.400 2649.440 23.470 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 624.750 197.100 625.070 197.160 ;
        RECT 2663.470 197.100 2663.790 197.160 ;
        RECT 624.750 196.960 2663.790 197.100 ;
        RECT 624.750 196.900 625.070 196.960 ;
        RECT 2663.470 196.900 2663.790 196.960 ;
      LAYER via ;
        RECT 624.780 196.900 625.040 197.160 ;
        RECT 2663.500 196.900 2663.760 197.160 ;
      LAYER met2 ;
        RECT 625.030 500.000 625.310 504.000 ;
        RECT 625.070 498.340 625.210 500.000 ;
        RECT 624.840 498.200 625.210 498.340 ;
        RECT 624.840 197.190 624.980 498.200 ;
        RECT 624.780 196.870 625.040 197.190 ;
        RECT 2663.500 196.870 2663.760 197.190 ;
        RECT 2663.560 82.870 2663.700 196.870 ;
        RECT 2663.560 82.730 2666.000 82.870 ;
        RECT 2665.860 2.400 2666.000 82.730 ;
        RECT 2665.650 -4.800 2666.210 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 410.850 761.160 411.170 761.220 ;
        RECT 484.450 761.160 484.770 761.220 ;
        RECT 410.850 761.020 484.770 761.160 ;
        RECT 410.850 760.960 411.170 761.020 ;
        RECT 484.450 760.960 484.770 761.020 ;
        RECT 475.940 498.820 476.260 499.080 ;
        RECT 476.030 497.660 476.170 498.820 ;
        RECT 475.340 497.520 476.170 497.660 ;
        RECT 475.340 497.380 475.480 497.520 ;
        RECT 475.250 497.120 475.570 497.380 ;
        RECT 581.970 486.780 582.290 486.840 ;
        RECT 496.730 486.640 582.290 486.780 ;
        RECT 466.970 486.440 467.290 486.500 ;
        RECT 475.250 486.440 475.570 486.500 ;
        RECT 496.730 486.440 496.870 486.640 ;
        RECT 581.970 486.580 582.290 486.640 ;
        RECT 466.970 486.300 496.870 486.440 ;
        RECT 466.970 486.240 467.290 486.300 ;
        RECT 475.250 486.240 475.570 486.300 ;
        RECT 410.850 484.740 411.170 484.800 ;
        RECT 410.850 484.600 433.620 484.740 ;
        RECT 410.850 484.540 411.170 484.600 ;
        RECT 433.480 484.060 433.620 484.600 ;
        RECT 466.970 484.060 467.290 484.120 ;
        RECT 433.480 483.920 467.290 484.060 ;
        RECT 466.970 483.860 467.290 483.920 ;
        RECT 581.970 482.700 582.290 482.760 ;
        RECT 584.270 482.700 584.590 482.760 ;
        RECT 581.970 482.560 584.590 482.700 ;
        RECT 581.970 482.500 582.290 482.560 ;
        RECT 584.270 482.500 584.590 482.560 ;
        RECT 584.270 461.280 584.590 461.340 ;
        RECT 876.370 461.280 876.690 461.340 ;
        RECT 584.270 461.140 876.690 461.280 ;
        RECT 584.270 461.080 584.590 461.140 ;
        RECT 876.370 461.080 876.690 461.140 ;
      LAYER via ;
        RECT 410.880 760.960 411.140 761.220 ;
        RECT 484.480 760.960 484.740 761.220 ;
        RECT 475.970 498.820 476.230 499.080 ;
        RECT 475.280 497.120 475.540 497.380 ;
        RECT 467.000 486.240 467.260 486.500 ;
        RECT 475.280 486.240 475.540 486.500 ;
        RECT 582.000 486.580 582.260 486.840 ;
        RECT 410.880 484.540 411.140 484.800 ;
        RECT 467.000 483.860 467.260 484.120 ;
        RECT 582.000 482.500 582.260 482.760 ;
        RECT 584.300 482.500 584.560 482.760 ;
        RECT 584.300 461.080 584.560 461.340 ;
        RECT 876.400 461.080 876.660 461.340 ;
      LAYER met2 ;
        RECT 410.880 760.930 411.140 761.250 ;
        RECT 484.480 760.930 484.740 761.250 ;
        RECT 410.940 484.830 411.080 760.930 ;
        RECT 484.540 749.770 484.680 760.930 ;
        RECT 485.190 749.770 485.470 750.000 ;
        RECT 484.540 749.630 485.470 749.770 ;
        RECT 485.190 746.000 485.470 749.630 ;
        RECT 475.990 500.000 476.270 504.000 ;
        RECT 476.030 499.110 476.170 500.000 ;
        RECT 475.970 498.790 476.230 499.110 ;
        RECT 475.280 497.090 475.540 497.410 ;
        RECT 475.340 486.530 475.480 497.090 ;
        RECT 582.000 486.550 582.260 486.870 ;
        RECT 467.000 486.210 467.260 486.530 ;
        RECT 475.280 486.210 475.540 486.530 ;
        RECT 410.880 484.510 411.140 484.830 ;
        RECT 467.060 484.150 467.200 486.210 ;
        RECT 467.000 483.830 467.260 484.150 ;
        RECT 582.060 482.790 582.200 486.550 ;
        RECT 582.000 482.470 582.260 482.790 ;
        RECT 584.300 482.470 584.560 482.790 ;
        RECT 584.360 461.370 584.500 482.470 ;
        RECT 584.300 461.050 584.560 461.370 ;
        RECT 876.400 461.050 876.660 461.370 ;
        RECT 876.460 17.410 876.600 461.050 ;
        RECT 876.460 17.270 877.520 17.410 ;
        RECT 877.380 2.400 877.520 17.270 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.410 500.000 626.690 504.000 ;
        RECT 626.450 499.645 626.590 500.000 ;
        RECT 626.380 499.275 626.660 499.645 ;
        RECT 2677.290 396.595 2677.570 396.965 ;
        RECT 2677.360 82.870 2677.500 396.595 ;
        RECT 2677.360 82.730 2682.560 82.870 ;
        RECT 2682.420 2.400 2682.560 82.730 ;
        RECT 2682.210 -4.800 2682.770 2.400 ;
      LAYER via2 ;
        RECT 626.380 499.320 626.660 499.600 ;
        RECT 2677.290 396.640 2677.570 396.920 ;
      LAYER met3 ;
        RECT 624.030 499.610 624.410 499.620 ;
        RECT 626.355 499.610 626.685 499.625 ;
        RECT 624.030 499.310 626.685 499.610 ;
        RECT 624.030 499.300 624.410 499.310 ;
        RECT 626.355 499.295 626.685 499.310 ;
        RECT 624.030 396.930 624.410 396.940 ;
        RECT 2677.265 396.930 2677.595 396.945 ;
        RECT 624.030 396.630 2677.595 396.930 ;
        RECT 624.030 396.620 624.410 396.630 ;
        RECT 2677.265 396.615 2677.595 396.630 ;
      LAYER via3 ;
        RECT 624.060 499.300 624.380 499.620 ;
        RECT 624.060 396.620 624.380 396.940 ;
      LAYER met4 ;
        RECT 624.055 499.295 624.385 499.625 ;
        RECT 624.070 396.945 624.370 499.295 ;
        RECT 624.055 396.615 624.385 396.945 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.740 499.500 628.060 499.760 ;
        RECT 627.830 499.360 627.970 499.500 ;
        RECT 627.830 499.220 628.660 499.360 ;
        RECT 628.520 497.040 628.660 499.220 ;
        RECT 628.430 496.780 628.750 497.040 ;
        RECT 628.430 31.520 628.750 31.580 ;
        RECT 2698.890 31.520 2699.210 31.580 ;
        RECT 628.430 31.380 2699.210 31.520 ;
        RECT 628.430 31.320 628.750 31.380 ;
        RECT 2698.890 31.320 2699.210 31.380 ;
      LAYER via ;
        RECT 627.770 499.500 628.030 499.760 ;
        RECT 628.460 496.780 628.720 497.040 ;
        RECT 628.460 31.320 628.720 31.580 ;
        RECT 2698.920 31.320 2699.180 31.580 ;
      LAYER met2 ;
        RECT 627.790 500.000 628.070 504.000 ;
        RECT 627.830 499.790 627.970 500.000 ;
        RECT 627.770 499.470 628.030 499.790 ;
        RECT 628.460 496.750 628.720 497.070 ;
        RECT 628.520 31.610 628.660 496.750 ;
        RECT 628.460 31.290 628.720 31.610 ;
        RECT 2698.920 31.290 2699.180 31.610 ;
        RECT 2698.980 2.400 2699.120 31.290 ;
        RECT 2698.770 -4.800 2699.330 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.120 498.820 629.440 499.080 ;
        RECT 629.210 497.660 629.350 498.820 ;
        RECT 631.190 497.660 631.510 497.720 ;
        RECT 629.210 497.520 631.510 497.660 ;
        RECT 631.190 497.460 631.510 497.520 ;
        RECT 631.190 196.760 631.510 196.820 ;
        RECT 2711.770 196.760 2712.090 196.820 ;
        RECT 631.190 196.620 2712.090 196.760 ;
        RECT 631.190 196.560 631.510 196.620 ;
        RECT 2711.770 196.560 2712.090 196.620 ;
      LAYER via ;
        RECT 629.150 498.820 629.410 499.080 ;
        RECT 631.220 497.460 631.480 497.720 ;
        RECT 631.220 196.560 631.480 196.820 ;
        RECT 2711.800 196.560 2712.060 196.820 ;
      LAYER met2 ;
        RECT 629.170 500.000 629.450 504.000 ;
        RECT 629.210 499.110 629.350 500.000 ;
        RECT 629.150 498.790 629.410 499.110 ;
        RECT 631.220 497.430 631.480 497.750 ;
        RECT 631.280 196.850 631.420 497.430 ;
        RECT 631.220 196.530 631.480 196.850 ;
        RECT 2711.800 196.530 2712.060 196.850 ;
        RECT 2711.860 82.870 2712.000 196.530 ;
        RECT 2711.860 82.730 2715.680 82.870 ;
        RECT 2715.540 2.400 2715.680 82.730 ;
        RECT 2715.330 -4.800 2715.890 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.730 496.980 631.050 497.040 ;
        RECT 632.110 496.980 632.430 497.040 ;
        RECT 630.730 496.840 632.430 496.980 ;
        RECT 630.730 496.780 631.050 496.840 ;
        RECT 632.110 496.780 632.430 496.840 ;
        RECT 632.110 438.500 632.430 438.560 ;
        RECT 2726.030 438.500 2726.350 438.560 ;
        RECT 632.110 438.360 2726.350 438.500 ;
        RECT 632.110 438.300 632.430 438.360 ;
        RECT 2726.030 438.300 2726.350 438.360 ;
        RECT 2726.030 17.920 2726.350 17.980 ;
        RECT 2732.010 17.920 2732.330 17.980 ;
        RECT 2726.030 17.780 2732.330 17.920 ;
        RECT 2726.030 17.720 2726.350 17.780 ;
        RECT 2732.010 17.720 2732.330 17.780 ;
      LAYER via ;
        RECT 630.760 496.780 631.020 497.040 ;
        RECT 632.140 496.780 632.400 497.040 ;
        RECT 632.140 438.300 632.400 438.560 ;
        RECT 2726.060 438.300 2726.320 438.560 ;
        RECT 2726.060 17.720 2726.320 17.980 ;
        RECT 2732.040 17.720 2732.300 17.980 ;
      LAYER met2 ;
        RECT 630.550 500.000 630.830 504.000 ;
        RECT 630.590 498.340 630.730 500.000 ;
        RECT 630.590 498.200 630.960 498.340 ;
        RECT 630.820 497.070 630.960 498.200 ;
        RECT 630.760 496.750 631.020 497.070 ;
        RECT 632.140 496.750 632.400 497.070 ;
        RECT 632.200 438.590 632.340 496.750 ;
        RECT 632.140 438.270 632.400 438.590 ;
        RECT 2726.060 438.270 2726.320 438.590 ;
        RECT 2726.120 18.010 2726.260 438.270 ;
        RECT 2726.060 17.690 2726.320 18.010 ;
        RECT 2732.040 17.690 2732.300 18.010 ;
        RECT 2732.100 2.400 2732.240 17.690 ;
        RECT 2731.890 -4.800 2732.450 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 631.880 499.500 632.200 499.760 ;
        RECT 631.970 499.020 632.110 499.500 ;
        RECT 631.970 498.880 633.030 499.020 ;
        RECT 632.110 498.000 632.430 498.060 ;
        RECT 632.890 498.000 633.030 498.880 ;
        RECT 632.110 497.860 633.030 498.000 ;
        RECT 632.110 497.800 632.430 497.860 ;
        RECT 631.650 438.160 631.970 438.220 ;
        RECT 2746.270 438.160 2746.590 438.220 ;
        RECT 631.650 438.020 2746.590 438.160 ;
        RECT 631.650 437.960 631.970 438.020 ;
        RECT 2746.270 437.960 2746.590 438.020 ;
      LAYER via ;
        RECT 631.910 499.500 632.170 499.760 ;
        RECT 632.140 497.800 632.400 498.060 ;
        RECT 631.680 437.960 631.940 438.220 ;
        RECT 2746.300 437.960 2746.560 438.220 ;
      LAYER met2 ;
        RECT 631.930 500.000 632.210 504.000 ;
        RECT 631.970 499.790 632.110 500.000 ;
        RECT 631.910 499.470 632.170 499.790 ;
        RECT 632.140 497.770 632.400 498.090 ;
        RECT 632.200 497.490 632.340 497.770 ;
        RECT 631.740 497.350 632.340 497.490 ;
        RECT 631.740 438.250 631.880 497.350 ;
        RECT 631.680 437.930 631.940 438.250 ;
        RECT 2746.300 437.930 2746.560 438.250 ;
        RECT 2746.360 82.870 2746.500 437.930 ;
        RECT 2746.360 82.730 2748.800 82.870 ;
        RECT 2748.660 2.400 2748.800 82.730 ;
        RECT 2748.450 -4.800 2749.010 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.310 500.000 633.590 504.000 ;
        RECT 633.350 499.815 633.490 500.000 ;
        RECT 633.280 499.445 633.560 499.815 ;
        RECT 2760.090 195.995 2760.370 196.365 ;
        RECT 2760.160 82.870 2760.300 195.995 ;
        RECT 2760.160 82.730 2765.360 82.870 ;
        RECT 2765.220 2.400 2765.360 82.730 ;
        RECT 2765.010 -4.800 2765.570 2.400 ;
      LAYER via2 ;
        RECT 633.280 499.490 633.560 499.770 ;
        RECT 2760.090 196.040 2760.370 196.320 ;
      LAYER met3 ;
        RECT 633.255 499.620 633.585 499.795 ;
        RECT 633.230 499.610 633.610 499.620 ;
        RECT 633.230 499.310 633.870 499.610 ;
        RECT 633.230 499.300 633.610 499.310 ;
        RECT 631.390 196.330 631.770 196.340 ;
        RECT 2760.065 196.330 2760.395 196.345 ;
        RECT 631.390 196.030 2760.395 196.330 ;
        RECT 631.390 196.020 631.770 196.030 ;
        RECT 2760.065 196.015 2760.395 196.030 ;
      LAYER via3 ;
        RECT 633.260 499.300 633.580 499.620 ;
        RECT 631.420 196.020 631.740 196.340 ;
      LAYER met4 ;
        RECT 633.255 499.295 633.585 499.625 ;
        RECT 633.270 494.850 633.570 499.295 ;
        RECT 631.430 494.550 633.570 494.850 ;
        RECT 631.430 196.345 631.730 494.550 ;
        RECT 631.415 196.015 631.745 196.345 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.730 499.900 636.940 500.040 ;
        RECT 634.730 499.760 634.870 499.900 ;
        RECT 634.640 499.500 634.960 499.760 ;
        RECT 636.800 499.360 636.940 499.900 ;
        RECT 638.090 499.360 638.410 499.420 ;
        RECT 636.800 499.220 638.410 499.360 ;
        RECT 638.090 499.160 638.410 499.220 ;
        RECT 638.090 31.180 638.410 31.240 ;
        RECT 2781.690 31.180 2782.010 31.240 ;
        RECT 638.090 31.040 2782.010 31.180 ;
        RECT 638.090 30.980 638.410 31.040 ;
        RECT 2781.690 30.980 2782.010 31.040 ;
      LAYER via ;
        RECT 634.670 499.500 634.930 499.760 ;
        RECT 638.120 499.160 638.380 499.420 ;
        RECT 638.120 30.980 638.380 31.240 ;
        RECT 2781.720 30.980 2781.980 31.240 ;
      LAYER met2 ;
        RECT 634.690 500.000 634.970 504.000 ;
        RECT 634.730 499.790 634.870 500.000 ;
        RECT 634.670 499.470 634.930 499.790 ;
        RECT 638.120 499.130 638.380 499.450 ;
        RECT 638.180 31.270 638.320 499.130 ;
        RECT 638.120 30.950 638.380 31.270 ;
        RECT 2781.720 30.950 2781.980 31.270 ;
        RECT 2781.780 2.400 2781.920 30.950 ;
        RECT 2781.570 -4.800 2782.130 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.020 499.500 636.340 499.760 ;
        RECT 636.110 498.060 636.250 499.500 ;
        RECT 636.110 497.860 636.570 498.060 ;
        RECT 636.250 497.800 636.570 497.860 ;
        RECT 636.250 444.620 636.570 444.680 ;
        RECT 637.630 444.620 637.950 444.680 ;
        RECT 636.250 444.480 637.950 444.620 ;
        RECT 636.250 444.420 636.570 444.480 ;
        RECT 637.630 444.420 637.950 444.480 ;
        RECT 637.630 30.840 637.950 30.900 ;
        RECT 2798.250 30.840 2798.570 30.900 ;
        RECT 637.630 30.700 2798.570 30.840 ;
        RECT 637.630 30.640 637.950 30.700 ;
        RECT 2798.250 30.640 2798.570 30.700 ;
      LAYER via ;
        RECT 636.050 499.500 636.310 499.760 ;
        RECT 636.280 497.800 636.540 498.060 ;
        RECT 636.280 444.420 636.540 444.680 ;
        RECT 637.660 444.420 637.920 444.680 ;
        RECT 637.660 30.640 637.920 30.900 ;
        RECT 2798.280 30.640 2798.540 30.900 ;
      LAYER met2 ;
        RECT 636.070 500.000 636.350 504.000 ;
        RECT 636.110 499.790 636.250 500.000 ;
        RECT 636.050 499.470 636.310 499.790 ;
        RECT 636.280 497.770 636.540 498.090 ;
        RECT 636.340 444.710 636.480 497.770 ;
        RECT 636.280 444.390 636.540 444.710 ;
        RECT 637.660 444.390 637.920 444.710 ;
        RECT 637.720 30.930 637.860 444.390 ;
        RECT 637.660 30.610 637.920 30.930 ;
        RECT 2798.280 30.610 2798.540 30.930 ;
        RECT 2798.340 2.400 2798.480 30.610 ;
        RECT 2798.130 -4.800 2798.690 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 411.310 759.120 411.630 759.180 ;
        RECT 490.890 759.120 491.210 759.180 ;
        RECT 411.310 758.980 491.210 759.120 ;
        RECT 411.310 758.920 411.630 758.980 ;
        RECT 490.890 758.920 491.210 758.980 ;
        RECT 476.630 483.040 476.950 483.100 ;
        RECT 448.430 482.900 476.950 483.040 ;
        RECT 411.310 482.700 411.630 482.760 ;
        RECT 448.430 482.700 448.570 482.900 ;
        RECT 476.630 482.840 476.950 482.900 ;
        RECT 411.310 482.560 448.570 482.700 ;
        RECT 411.310 482.500 411.630 482.560 ;
        RECT 476.630 476.240 476.950 476.300 ;
        RECT 480.770 476.240 481.090 476.300 ;
        RECT 476.630 476.100 481.090 476.240 ;
        RECT 476.630 476.040 476.950 476.100 ;
        RECT 480.770 476.040 481.090 476.100 ;
        RECT 480.770 447.680 481.090 447.740 ;
        RECT 890.170 447.680 890.490 447.740 ;
        RECT 480.770 447.540 890.490 447.680 ;
        RECT 480.770 447.480 481.090 447.540 ;
        RECT 890.170 447.480 890.490 447.540 ;
      LAYER via ;
        RECT 411.340 758.920 411.600 759.180 ;
        RECT 490.920 758.920 491.180 759.180 ;
        RECT 411.340 482.500 411.600 482.760 ;
        RECT 476.660 482.840 476.920 483.100 ;
        RECT 476.660 476.040 476.920 476.300 ;
        RECT 480.800 476.040 481.060 476.300 ;
        RECT 480.800 447.480 481.060 447.740 ;
        RECT 890.200 447.480 890.460 447.740 ;
      LAYER met2 ;
        RECT 411.340 758.890 411.600 759.210 ;
        RECT 490.920 758.890 491.180 759.210 ;
        RECT 411.400 482.790 411.540 758.890 ;
        RECT 490.980 750.000 491.120 758.890 ;
        RECT 490.710 749.630 491.120 750.000 ;
        RECT 490.710 746.000 490.990 749.630 ;
        RECT 477.370 500.000 477.650 504.000 ;
        RECT 477.410 499.645 477.550 500.000 ;
        RECT 477.340 499.275 477.620 499.645 ;
        RECT 476.650 491.115 476.930 491.485 ;
        RECT 476.720 483.130 476.860 491.115 ;
        RECT 476.660 482.810 476.920 483.130 ;
        RECT 411.340 482.470 411.600 482.790 ;
        RECT 476.720 476.330 476.860 482.810 ;
        RECT 476.660 476.010 476.920 476.330 ;
        RECT 480.800 476.010 481.060 476.330 ;
        RECT 480.860 447.770 481.000 476.010 ;
        RECT 480.800 447.450 481.060 447.770 ;
        RECT 890.200 447.450 890.460 447.770 ;
        RECT 890.260 82.870 890.400 447.450 ;
        RECT 890.260 82.730 894.080 82.870 ;
        RECT 893.940 2.400 894.080 82.730 ;
        RECT 893.730 -4.800 894.290 2.400 ;
      LAYER via2 ;
        RECT 477.340 499.320 477.620 499.600 ;
        RECT 476.650 491.160 476.930 491.440 ;
      LAYER met3 ;
        RECT 475.910 499.610 476.290 499.620 ;
        RECT 477.315 499.610 477.645 499.625 ;
        RECT 475.910 499.310 477.645 499.610 ;
        RECT 475.910 499.300 476.290 499.310 ;
        RECT 477.315 499.295 477.645 499.310 ;
        RECT 475.910 491.450 476.290 491.460 ;
        RECT 476.625 491.450 476.955 491.465 ;
        RECT 475.910 491.150 476.955 491.450 ;
        RECT 475.910 491.140 476.290 491.150 ;
        RECT 476.625 491.135 476.955 491.150 ;
      LAYER via3 ;
        RECT 475.940 499.300 476.260 499.620 ;
        RECT 475.940 491.140 476.260 491.460 ;
      LAYER met4 ;
        RECT 475.935 499.295 476.265 499.625 ;
        RECT 475.950 491.465 476.250 499.295 ;
        RECT 475.935 491.135 476.265 491.465 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.550 760.820 408.870 760.880 ;
        RECT 495.490 760.820 495.810 760.880 ;
        RECT 408.550 760.680 495.810 760.820 ;
        RECT 408.550 760.620 408.870 760.680 ;
        RECT 495.490 760.620 495.810 760.680 ;
        RECT 478.700 499.500 479.020 499.760 ;
        RECT 408.550 496.300 408.870 496.360 ;
        RECT 478.790 496.300 478.930 499.500 ;
        RECT 480.310 496.300 480.630 496.360 ;
        RECT 408.550 496.160 480.630 496.300 ;
        RECT 408.550 496.100 408.870 496.160 ;
        RECT 480.310 496.100 480.630 496.160 ;
        RECT 479.390 472.840 479.710 472.900 ;
        RECT 480.310 472.840 480.630 472.900 ;
        RECT 479.390 472.700 480.630 472.840 ;
        RECT 479.390 472.640 479.710 472.700 ;
        RECT 480.310 472.640 480.630 472.700 ;
        RECT 479.390 447.340 479.710 447.400 ;
        RECT 903.970 447.340 904.290 447.400 ;
        RECT 479.390 447.200 904.290 447.340 ;
        RECT 479.390 447.140 479.710 447.200 ;
        RECT 903.970 447.140 904.290 447.200 ;
        RECT 903.970 16.900 904.290 16.960 ;
        RECT 910.410 16.900 910.730 16.960 ;
        RECT 903.970 16.760 910.730 16.900 ;
        RECT 903.970 16.700 904.290 16.760 ;
        RECT 910.410 16.700 910.730 16.760 ;
      LAYER via ;
        RECT 408.580 760.620 408.840 760.880 ;
        RECT 495.520 760.620 495.780 760.880 ;
        RECT 478.730 499.500 478.990 499.760 ;
        RECT 408.580 496.100 408.840 496.360 ;
        RECT 480.340 496.100 480.600 496.360 ;
        RECT 479.420 472.640 479.680 472.900 ;
        RECT 480.340 472.640 480.600 472.900 ;
        RECT 479.420 447.140 479.680 447.400 ;
        RECT 904.000 447.140 904.260 447.400 ;
        RECT 904.000 16.700 904.260 16.960 ;
        RECT 910.440 16.700 910.700 16.960 ;
      LAYER met2 ;
        RECT 408.580 760.590 408.840 760.910 ;
        RECT 495.520 760.590 495.780 760.910 ;
        RECT 408.640 545.090 408.780 760.590 ;
        RECT 495.580 749.770 495.720 760.590 ;
        RECT 496.230 749.770 496.510 750.000 ;
        RECT 495.580 749.630 496.510 749.770 ;
        RECT 496.230 746.000 496.510 749.630 ;
        RECT 408.180 544.950 408.780 545.090 ;
        RECT 408.180 531.370 408.320 544.950 ;
        RECT 408.180 531.230 408.780 531.370 ;
        RECT 408.640 496.390 408.780 531.230 ;
        RECT 478.750 500.000 479.030 504.000 ;
        RECT 478.790 499.790 478.930 500.000 ;
        RECT 478.730 499.470 478.990 499.790 ;
        RECT 408.580 496.070 408.840 496.390 ;
        RECT 480.340 496.070 480.600 496.390 ;
        RECT 480.400 472.930 480.540 496.070 ;
        RECT 479.420 472.610 479.680 472.930 ;
        RECT 480.340 472.610 480.600 472.930 ;
        RECT 479.480 447.430 479.620 472.610 ;
        RECT 479.420 447.110 479.680 447.430 ;
        RECT 904.000 447.110 904.260 447.430 ;
        RECT 904.060 16.990 904.200 447.110 ;
        RECT 904.000 16.670 904.260 16.990 ;
        RECT 910.440 16.670 910.700 16.990 ;
        RECT 910.500 2.400 910.640 16.670 ;
        RECT 910.290 -4.800 910.850 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 760.480 407.490 760.540 ;
        RECT 501.010 760.480 501.330 760.540 ;
        RECT 407.170 760.340 501.330 760.480 ;
        RECT 407.170 760.280 407.490 760.340 ;
        RECT 501.010 760.280 501.330 760.340 ;
        RECT 407.170 499.700 407.490 499.760 ;
        RECT 411.770 499.700 412.090 499.760 ;
        RECT 407.170 499.560 412.090 499.700 ;
        RECT 407.170 499.500 407.490 499.560 ;
        RECT 411.770 499.500 412.090 499.560 ;
        RECT 480.080 499.500 480.400 499.760 ;
        RECT 480.170 499.080 480.310 499.500 ;
        RECT 479.850 498.880 480.310 499.080 ;
        RECT 479.850 498.820 480.170 498.880 ;
        RECT 411.770 481.000 412.090 481.060 ;
        RECT 479.850 481.000 480.170 481.060 ;
        RECT 411.770 480.860 480.170 481.000 ;
        RECT 411.770 480.800 412.090 480.860 ;
        RECT 479.850 480.800 480.170 480.860 ;
        RECT 480.310 32.540 480.630 32.600 ;
        RECT 926.970 32.540 927.290 32.600 ;
        RECT 480.310 32.400 927.290 32.540 ;
        RECT 480.310 32.340 480.630 32.400 ;
        RECT 926.970 32.340 927.290 32.400 ;
      LAYER via ;
        RECT 407.200 760.280 407.460 760.540 ;
        RECT 501.040 760.280 501.300 760.540 ;
        RECT 407.200 499.500 407.460 499.760 ;
        RECT 411.800 499.500 412.060 499.760 ;
        RECT 480.110 499.500 480.370 499.760 ;
        RECT 479.880 498.820 480.140 499.080 ;
        RECT 411.800 480.800 412.060 481.060 ;
        RECT 479.880 480.800 480.140 481.060 ;
        RECT 480.340 32.340 480.600 32.600 ;
        RECT 927.000 32.340 927.260 32.600 ;
      LAYER met2 ;
        RECT 407.200 760.250 407.460 760.570 ;
        RECT 501.040 760.250 501.300 760.570 ;
        RECT 407.260 565.870 407.400 760.250 ;
        RECT 501.100 749.770 501.240 760.250 ;
        RECT 501.750 749.770 502.030 750.000 ;
        RECT 501.100 749.630 502.030 749.770 ;
        RECT 501.750 746.000 502.030 749.630 ;
        RECT 407.260 565.730 407.860 565.870 ;
        RECT 407.720 545.170 407.860 565.730 ;
        RECT 407.260 545.030 407.860 545.170 ;
        RECT 407.260 499.790 407.400 545.030 ;
        RECT 480.130 500.000 480.410 504.000 ;
        RECT 480.170 499.790 480.310 500.000 ;
        RECT 407.200 499.470 407.460 499.790 ;
        RECT 411.800 499.470 412.060 499.790 ;
        RECT 480.110 499.470 480.370 499.790 ;
        RECT 411.860 481.090 412.000 499.470 ;
        RECT 479.880 498.790 480.140 499.110 ;
        RECT 479.940 481.090 480.080 498.790 ;
        RECT 411.800 480.770 412.060 481.090 ;
        RECT 479.880 480.770 480.140 481.090 ;
        RECT 479.940 472.330 480.080 480.770 ;
        RECT 479.940 472.190 480.540 472.330 ;
        RECT 480.400 32.630 480.540 472.190 ;
        RECT 480.340 32.310 480.600 32.630 ;
        RECT 927.000 32.310 927.260 32.630 ;
        RECT 927.060 2.400 927.200 32.310 ;
        RECT 926.850 -4.800 927.410 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 411.770 761.500 412.090 761.560 ;
        RECT 506.530 761.500 506.850 761.560 ;
        RECT 411.770 761.360 506.850 761.500 ;
        RECT 411.770 761.300 412.090 761.360 ;
        RECT 506.530 761.300 506.850 761.360 ;
        RECT 409.470 507.520 409.790 507.580 ;
        RECT 411.770 507.520 412.090 507.580 ;
        RECT 409.470 507.380 412.090 507.520 ;
        RECT 409.470 507.320 409.790 507.380 ;
        RECT 411.770 507.320 412.090 507.380 ;
        RECT 481.460 499.500 481.780 499.760 ;
        RECT 407.170 499.020 407.490 499.080 ;
        RECT 409.470 499.020 409.790 499.080 ;
        RECT 407.170 498.880 409.790 499.020 ;
        RECT 407.170 498.820 407.490 498.880 ;
        RECT 409.470 498.820 409.790 498.880 ;
        RECT 481.550 497.660 481.690 499.500 ;
        RECT 482.150 497.660 482.470 497.720 ;
        RECT 481.550 497.520 482.470 497.660 ;
        RECT 482.150 497.460 482.470 497.520 ;
        RECT 407.170 481.340 407.490 481.400 ;
        RECT 482.150 481.340 482.470 481.400 ;
        RECT 407.170 481.200 482.470 481.340 ;
        RECT 407.170 481.140 407.490 481.200 ;
        RECT 482.150 481.140 482.470 481.200 ;
        RECT 479.850 471.820 480.170 471.880 ;
        RECT 482.610 471.820 482.930 471.880 ;
        RECT 479.850 471.680 482.930 471.820 ;
        RECT 479.850 471.620 480.170 471.680 ;
        RECT 482.610 471.620 482.930 471.680 ;
        RECT 479.850 32.200 480.170 32.260 ;
        RECT 943.530 32.200 943.850 32.260 ;
        RECT 479.850 32.060 943.850 32.200 ;
        RECT 479.850 32.000 480.170 32.060 ;
        RECT 943.530 32.000 943.850 32.060 ;
      LAYER via ;
        RECT 411.800 761.300 412.060 761.560 ;
        RECT 506.560 761.300 506.820 761.560 ;
        RECT 409.500 507.320 409.760 507.580 ;
        RECT 411.800 507.320 412.060 507.580 ;
        RECT 481.490 499.500 481.750 499.760 ;
        RECT 407.200 498.820 407.460 499.080 ;
        RECT 409.500 498.820 409.760 499.080 ;
        RECT 482.180 497.460 482.440 497.720 ;
        RECT 407.200 481.140 407.460 481.400 ;
        RECT 482.180 481.140 482.440 481.400 ;
        RECT 479.880 471.620 480.140 471.880 ;
        RECT 482.640 471.620 482.900 471.880 ;
        RECT 479.880 32.000 480.140 32.260 ;
        RECT 943.560 32.000 943.820 32.260 ;
      LAYER met2 ;
        RECT 411.800 761.270 412.060 761.590 ;
        RECT 506.560 761.270 506.820 761.590 ;
        RECT 411.860 507.610 412.000 761.270 ;
        RECT 506.620 749.770 506.760 761.270 ;
        RECT 507.270 749.770 507.550 750.000 ;
        RECT 506.620 749.630 507.550 749.770 ;
        RECT 507.270 746.000 507.550 749.630 ;
        RECT 409.500 507.290 409.760 507.610 ;
        RECT 411.800 507.290 412.060 507.610 ;
        RECT 409.560 499.110 409.700 507.290 ;
        RECT 481.510 500.000 481.790 504.000 ;
        RECT 481.550 499.790 481.690 500.000 ;
        RECT 481.490 499.470 481.750 499.790 ;
        RECT 407.200 498.790 407.460 499.110 ;
        RECT 409.500 498.790 409.760 499.110 ;
        RECT 407.260 481.430 407.400 498.790 ;
        RECT 482.180 497.430 482.440 497.750 ;
        RECT 482.240 481.430 482.380 497.430 ;
        RECT 407.200 481.110 407.460 481.430 ;
        RECT 482.180 481.110 482.440 481.430 ;
        RECT 482.240 476.170 482.380 481.110 ;
        RECT 482.240 476.030 482.840 476.170 ;
        RECT 482.700 471.910 482.840 476.030 ;
        RECT 479.880 471.590 480.140 471.910 ;
        RECT 482.640 471.590 482.900 471.910 ;
        RECT 479.940 32.290 480.080 471.590 ;
        RECT 479.880 31.970 480.140 32.290 ;
        RECT 943.560 31.970 943.820 32.290 ;
        RECT 943.620 2.400 943.760 31.970 ;
        RECT 943.410 -4.800 943.970 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 482.840 499.700 483.160 499.760 ;
        RECT 482.840 499.560 483.760 499.700 ;
        RECT 482.840 499.500 483.160 499.560 ;
        RECT 483.620 498.400 483.760 499.560 ;
        RECT 483.530 498.140 483.850 498.400 ;
        RECT 483.530 479.300 483.850 479.360 ;
        RECT 485.830 479.300 486.150 479.360 ;
        RECT 483.530 479.160 486.150 479.300 ;
        RECT 483.530 479.100 483.850 479.160 ;
        RECT 485.830 479.100 486.150 479.160 ;
        RECT 485.830 460.940 486.150 461.000 ;
        RECT 625.210 460.940 625.530 461.000 ;
        RECT 485.830 460.800 625.530 460.940 ;
        RECT 485.830 460.740 486.150 460.800 ;
        RECT 625.210 460.740 625.530 460.800 ;
        RECT 625.210 455.500 625.530 455.560 ;
        RECT 959.170 455.500 959.490 455.560 ;
        RECT 625.210 455.360 959.490 455.500 ;
        RECT 625.210 455.300 625.530 455.360 ;
        RECT 959.170 455.300 959.490 455.360 ;
      LAYER via ;
        RECT 482.870 499.500 483.130 499.760 ;
        RECT 483.560 498.140 483.820 498.400 ;
        RECT 483.560 479.100 483.820 479.360 ;
        RECT 485.860 479.100 486.120 479.360 ;
        RECT 485.860 460.740 486.120 461.000 ;
        RECT 625.240 460.740 625.500 461.000 ;
        RECT 625.240 455.300 625.500 455.560 ;
        RECT 959.200 455.300 959.460 455.560 ;
      LAYER met2 ;
        RECT 513.450 761.075 513.730 761.445 ;
        RECT 512.790 749.770 513.070 750.000 ;
        RECT 513.520 749.770 513.660 761.075 ;
        RECT 512.790 749.630 513.660 749.770 ;
        RECT 512.790 746.000 513.070 749.630 ;
        RECT 482.890 500.000 483.170 504.000 ;
        RECT 482.930 499.790 483.070 500.000 ;
        RECT 482.870 499.470 483.130 499.790 ;
        RECT 483.560 498.110 483.820 498.430 ;
        RECT 483.620 479.390 483.760 498.110 ;
        RECT 483.560 479.070 483.820 479.390 ;
        RECT 485.860 479.070 486.120 479.390 ;
        RECT 485.920 461.030 486.060 479.070 ;
        RECT 625.230 461.875 625.510 462.245 ;
        RECT 625.300 461.030 625.440 461.875 ;
        RECT 485.860 460.710 486.120 461.030 ;
        RECT 625.240 460.710 625.500 461.030 ;
        RECT 625.300 455.590 625.440 460.710 ;
        RECT 625.240 455.270 625.500 455.590 ;
        RECT 959.200 455.270 959.460 455.590 ;
        RECT 959.260 17.410 959.400 455.270 ;
        RECT 959.260 17.270 960.320 17.410 ;
        RECT 960.180 2.400 960.320 17.270 ;
        RECT 959.970 -4.800 960.530 2.400 ;
      LAYER via2 ;
        RECT 513.450 761.120 513.730 761.400 ;
        RECT 625.230 461.920 625.510 462.200 ;
      LAYER met3 ;
        RECT 513.425 761.410 513.755 761.425 ;
        RECT 621.270 761.410 621.650 761.420 ;
        RECT 513.425 761.110 621.650 761.410 ;
        RECT 513.425 761.095 513.755 761.110 ;
        RECT 621.270 761.100 621.650 761.110 ;
        RECT 621.270 462.210 621.650 462.220 ;
        RECT 625.205 462.210 625.535 462.225 ;
        RECT 621.270 461.910 625.535 462.210 ;
        RECT 621.270 461.900 621.650 461.910 ;
        RECT 625.205 461.895 625.535 461.910 ;
      LAYER via3 ;
        RECT 621.300 761.100 621.620 761.420 ;
        RECT 621.300 461.900 621.620 462.220 ;
      LAYER met4 ;
        RECT 621.295 761.095 621.625 761.425 ;
        RECT 621.310 462.225 621.610 761.095 ;
        RECT 621.295 461.895 621.625 462.225 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.950 760.140 519.270 760.200 ;
        RECT 644.070 760.140 644.390 760.200 ;
        RECT 518.950 760.000 644.390 760.140 ;
        RECT 518.950 759.940 519.270 760.000 ;
        RECT 644.070 759.940 644.390 760.000 ;
        RECT 484.220 499.360 484.540 499.420 ;
        RECT 484.080 499.160 484.540 499.360 ;
        RECT 484.080 498.340 484.220 499.160 ;
        RECT 485.830 498.340 486.150 498.400 ;
        RECT 484.080 498.200 486.150 498.340 ;
        RECT 485.830 498.140 486.150 498.200 ;
        RECT 486.290 462.300 486.610 462.360 ;
        RECT 644.070 462.300 644.390 462.360 ;
        RECT 486.290 462.160 644.390 462.300 ;
        RECT 486.290 462.100 486.610 462.160 ;
        RECT 644.070 462.100 644.390 462.160 ;
        RECT 644.070 460.940 644.390 461.000 ;
        RECT 972.970 460.940 973.290 461.000 ;
        RECT 644.070 460.800 973.290 460.940 ;
        RECT 644.070 460.740 644.390 460.800 ;
        RECT 972.970 460.740 973.290 460.800 ;
      LAYER via ;
        RECT 518.980 759.940 519.240 760.200 ;
        RECT 644.100 759.940 644.360 760.200 ;
        RECT 484.250 499.160 484.510 499.420 ;
        RECT 485.860 498.140 486.120 498.400 ;
        RECT 486.320 462.100 486.580 462.360 ;
        RECT 644.100 462.100 644.360 462.360 ;
        RECT 644.100 460.740 644.360 461.000 ;
        RECT 973.000 460.740 973.260 461.000 ;
      LAYER met2 ;
        RECT 518.980 759.910 519.240 760.230 ;
        RECT 644.100 759.910 644.360 760.230 ;
        RECT 518.310 749.770 518.590 750.000 ;
        RECT 519.040 749.770 519.180 759.910 ;
        RECT 518.310 749.630 519.180 749.770 ;
        RECT 518.310 746.000 518.590 749.630 ;
        RECT 484.270 500.000 484.550 504.000 ;
        RECT 484.310 499.450 484.450 500.000 ;
        RECT 484.250 499.130 484.510 499.450 ;
        RECT 485.860 498.110 486.120 498.430 ;
        RECT 485.920 483.070 486.060 498.110 ;
        RECT 485.920 482.930 486.520 483.070 ;
        RECT 486.380 462.390 486.520 482.930 ;
        RECT 644.160 462.390 644.300 759.910 ;
        RECT 486.320 462.070 486.580 462.390 ;
        RECT 644.100 462.070 644.360 462.390 ;
        RECT 644.160 461.030 644.300 462.070 ;
        RECT 644.100 460.710 644.360 461.030 ;
        RECT 973.000 460.710 973.260 461.030 ;
        RECT 973.060 82.870 973.200 460.710 ;
        RECT 973.060 82.730 976.880 82.870 ;
        RECT 976.740 2.400 976.880 82.730 ;
        RECT 976.530 -4.800 977.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.010 760.480 524.330 760.540 ;
        RECT 641.770 760.480 642.090 760.540 ;
        RECT 524.010 760.340 642.090 760.480 ;
        RECT 524.010 760.280 524.330 760.340 ;
        RECT 641.770 760.280 642.090 760.340 ;
        RECT 485.600 499.360 485.920 499.420 ;
        RECT 485.460 499.160 485.920 499.360 ;
        RECT 485.460 498.740 485.600 499.160 ;
        RECT 485.370 498.480 485.690 498.740 ;
        RECT 485.370 427.620 485.690 427.680 ;
        RECT 641.770 427.620 642.090 427.680 ;
        RECT 485.370 427.480 662.470 427.620 ;
        RECT 485.370 427.420 485.690 427.480 ;
        RECT 641.770 427.420 642.090 427.480 ;
        RECT 662.330 426.260 662.470 427.480 ;
        RECT 986.770 426.260 987.090 426.320 ;
        RECT 662.330 426.120 987.090 426.260 ;
        RECT 986.770 426.060 987.090 426.120 ;
        RECT 986.770 16.900 987.090 16.960 ;
        RECT 993.210 16.900 993.530 16.960 ;
        RECT 986.770 16.760 993.530 16.900 ;
        RECT 986.770 16.700 987.090 16.760 ;
        RECT 993.210 16.700 993.530 16.760 ;
      LAYER via ;
        RECT 524.040 760.280 524.300 760.540 ;
        RECT 641.800 760.280 642.060 760.540 ;
        RECT 485.630 499.160 485.890 499.420 ;
        RECT 485.400 498.480 485.660 498.740 ;
        RECT 485.400 427.420 485.660 427.680 ;
        RECT 641.800 427.420 642.060 427.680 ;
        RECT 986.800 426.060 987.060 426.320 ;
        RECT 986.800 16.700 987.060 16.960 ;
        RECT 993.240 16.700 993.500 16.960 ;
      LAYER met2 ;
        RECT 524.040 760.250 524.300 760.570 ;
        RECT 641.800 760.250 642.060 760.570 ;
        RECT 524.100 750.000 524.240 760.250 ;
        RECT 523.830 749.630 524.240 750.000 ;
        RECT 523.830 746.000 524.110 749.630 ;
        RECT 485.650 500.000 485.930 504.000 ;
        RECT 485.690 499.450 485.830 500.000 ;
        RECT 485.630 499.130 485.890 499.450 ;
        RECT 485.400 498.450 485.660 498.770 ;
        RECT 485.460 427.710 485.600 498.450 ;
        RECT 641.860 449.210 642.000 760.250 ;
        RECT 641.400 449.070 642.000 449.210 ;
        RECT 641.400 446.490 641.540 449.070 ;
        RECT 641.400 446.350 642.000 446.490 ;
        RECT 641.860 427.710 642.000 446.350 ;
        RECT 485.400 427.390 485.660 427.710 ;
        RECT 641.800 427.390 642.060 427.710 ;
        RECT 986.800 426.030 987.060 426.350 ;
        RECT 986.860 16.990 987.000 426.030 ;
        RECT 986.800 16.670 987.060 16.990 ;
        RECT 993.240 16.670 993.500 16.990 ;
        RECT 993.300 2.400 993.440 16.670 ;
        RECT 993.090 -4.800 993.650 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.290 485.760 486.610 485.820 ;
        RECT 487.670 485.760 487.990 485.820 ;
        RECT 486.290 485.620 487.990 485.760 ;
        RECT 486.290 485.560 486.610 485.620 ;
        RECT 487.670 485.560 487.990 485.620 ;
        RECT 487.670 40.700 487.990 40.760 ;
        RECT 1009.770 40.700 1010.090 40.760 ;
        RECT 487.670 40.560 1010.090 40.700 ;
        RECT 487.670 40.500 487.990 40.560 ;
        RECT 1009.770 40.500 1010.090 40.560 ;
      LAYER via ;
        RECT 486.320 485.560 486.580 485.820 ;
        RECT 487.700 485.560 487.960 485.820 ;
        RECT 487.700 40.500 487.960 40.760 ;
        RECT 1009.800 40.500 1010.060 40.760 ;
      LAYER met2 ;
        RECT 528.630 759.035 528.910 759.405 ;
        RECT 528.700 749.770 528.840 759.035 ;
        RECT 529.350 749.770 529.630 750.000 ;
        RECT 528.700 749.630 529.630 749.770 ;
        RECT 529.350 746.000 529.630 749.630 ;
        RECT 487.030 500.000 487.310 504.000 ;
        RECT 487.070 499.815 487.210 500.000 ;
        RECT 487.000 499.445 487.280 499.815 ;
        RECT 486.770 498.850 487.050 498.965 ;
        RECT 486.380 498.710 487.050 498.850 ;
        RECT 486.380 485.850 486.520 498.710 ;
        RECT 486.770 498.595 487.050 498.710 ;
        RECT 486.320 485.530 486.580 485.850 ;
        RECT 487.700 485.530 487.960 485.850 ;
        RECT 487.760 481.965 487.900 485.530 ;
        RECT 487.690 481.595 487.970 481.965 ;
        RECT 487.760 40.790 487.900 481.595 ;
        RECT 487.700 40.470 487.960 40.790 ;
        RECT 1009.800 40.470 1010.060 40.790 ;
        RECT 1009.860 2.400 1010.000 40.470 ;
        RECT 1009.650 -4.800 1010.210 2.400 ;
      LAYER via2 ;
        RECT 528.630 759.080 528.910 759.360 ;
        RECT 487.000 499.490 487.280 499.770 ;
        RECT 486.770 498.640 487.050 498.920 ;
        RECT 487.690 481.640 487.970 481.920 ;
      LAYER met3 ;
        RECT 412.430 759.370 412.810 759.380 ;
        RECT 528.605 759.370 528.935 759.385 ;
        RECT 412.430 759.070 528.935 759.370 ;
        RECT 412.430 759.060 412.810 759.070 ;
        RECT 528.605 759.055 528.935 759.070 ;
        RECT 486.975 499.465 487.305 499.795 ;
        RECT 486.990 498.945 487.290 499.465 ;
        RECT 486.745 498.630 487.290 498.945 ;
        RECT 486.745 498.615 487.075 498.630 ;
        RECT 412.430 481.930 412.810 481.940 ;
        RECT 487.665 481.930 487.995 481.945 ;
        RECT 412.430 481.630 487.995 481.930 ;
        RECT 412.430 481.620 412.810 481.630 ;
        RECT 487.665 481.615 487.995 481.630 ;
      LAYER via3 ;
        RECT 412.460 759.060 412.780 759.380 ;
        RECT 412.460 481.620 412.780 481.940 ;
      LAYER met4 ;
        RECT 412.455 759.055 412.785 759.385 ;
        RECT 412.470 481.945 412.770 759.055 ;
        RECT 412.455 481.615 412.785 481.945 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 409.930 747.560 410.250 747.620 ;
        RECT 429.250 747.560 429.570 747.620 ;
        RECT 409.930 747.420 429.570 747.560 ;
        RECT 409.930 747.360 410.250 747.420 ;
        RECT 429.250 747.360 429.570 747.420 ;
        RECT 462.140 499.360 462.460 499.420 ;
        RECT 462.140 499.160 462.600 499.360 ;
        RECT 462.460 498.060 462.600 499.160 ;
        RECT 462.370 497.800 462.690 498.060 ;
        RECT 409.930 488.820 410.250 488.880 ;
        RECT 409.930 488.680 427.870 488.820 ;
        RECT 409.930 488.620 410.250 488.680 ;
        RECT 427.730 487.800 427.870 488.680 ;
        RECT 462.370 487.800 462.690 487.860 ;
        RECT 427.730 487.660 462.690 487.800 ;
        RECT 462.370 487.600 462.690 487.660 ;
        RECT 462.370 483.380 462.690 483.440 ;
        RECT 466.970 483.380 467.290 483.440 ;
        RECT 462.370 483.240 467.290 483.380 ;
        RECT 462.370 483.180 462.690 483.240 ;
        RECT 466.970 483.180 467.290 483.240 ;
        RECT 466.970 461.960 467.290 462.020 ;
        RECT 710.770 461.960 711.090 462.020 ;
        RECT 466.970 461.820 711.090 461.960 ;
        RECT 466.970 461.760 467.290 461.820 ;
        RECT 710.770 461.760 711.090 461.820 ;
      LAYER via ;
        RECT 409.960 747.360 410.220 747.620 ;
        RECT 429.280 747.360 429.540 747.620 ;
        RECT 462.170 499.160 462.430 499.420 ;
        RECT 462.400 497.800 462.660 498.060 ;
        RECT 409.960 488.620 410.220 488.880 ;
        RECT 462.400 487.600 462.660 487.860 ;
        RECT 462.400 483.180 462.660 483.440 ;
        RECT 467.000 483.180 467.260 483.440 ;
        RECT 467.000 461.760 467.260 462.020 ;
        RECT 710.800 461.760 711.060 462.020 ;
      LAYER met2 ;
        RECT 429.990 747.730 430.270 750.000 ;
        RECT 429.340 747.650 430.270 747.730 ;
        RECT 409.960 747.330 410.220 747.650 ;
        RECT 429.280 747.590 430.270 747.650 ;
        RECT 429.280 747.330 429.540 747.590 ;
        RECT 410.020 488.910 410.160 747.330 ;
        RECT 429.990 746.000 430.270 747.590 ;
        RECT 462.190 500.000 462.470 504.000 ;
        RECT 462.230 499.450 462.370 500.000 ;
        RECT 462.170 499.130 462.430 499.450 ;
        RECT 462.400 497.770 462.660 498.090 ;
        RECT 409.960 488.590 410.220 488.910 ;
        RECT 462.460 487.890 462.600 497.770 ;
        RECT 462.400 487.570 462.660 487.890 ;
        RECT 462.460 483.470 462.600 487.570 ;
        RECT 462.400 483.150 462.660 483.470 ;
        RECT 467.000 483.150 467.260 483.470 ;
        RECT 467.060 462.050 467.200 483.150 ;
        RECT 467.000 461.730 467.260 462.050 ;
        RECT 710.800 461.730 711.060 462.050 ;
        RECT 710.860 17.410 711.000 461.730 ;
        RECT 710.860 17.270 711.920 17.410 ;
        RECT 711.780 2.400 711.920 17.270 ;
        RECT 711.570 -4.800 712.130 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 488.360 499.700 488.680 499.760 ;
        RECT 488.360 499.560 489.510 499.700 ;
        RECT 488.360 499.500 488.680 499.560 ;
        RECT 489.370 497.720 489.510 499.560 ;
        RECT 489.370 497.520 489.830 497.720 ;
        RECT 489.510 497.460 489.830 497.520 ;
        RECT 483.070 474.200 483.390 474.260 ;
        RECT 489.510 474.200 489.830 474.260 ;
        RECT 483.070 474.060 489.830 474.200 ;
        RECT 483.070 474.000 483.390 474.060 ;
        RECT 489.510 474.000 489.830 474.060 ;
        RECT 483.070 40.360 483.390 40.420 ;
        RECT 1026.330 40.360 1026.650 40.420 ;
        RECT 483.070 40.220 1026.650 40.360 ;
        RECT 483.070 40.160 483.390 40.220 ;
        RECT 1026.330 40.160 1026.650 40.220 ;
      LAYER via ;
        RECT 488.390 499.500 488.650 499.760 ;
        RECT 489.540 497.460 489.800 497.720 ;
        RECT 483.100 474.000 483.360 474.260 ;
        RECT 489.540 474.000 489.800 474.260 ;
        RECT 483.100 40.160 483.360 40.420 ;
        RECT 1026.360 40.160 1026.620 40.420 ;
      LAYER met2 ;
        RECT 534.150 759.715 534.430 760.085 ;
        RECT 534.220 749.770 534.360 759.715 ;
        RECT 534.870 749.770 535.150 750.000 ;
        RECT 534.220 749.630 535.150 749.770 ;
        RECT 534.870 746.000 535.150 749.630 ;
        RECT 488.410 500.000 488.690 504.000 ;
        RECT 488.450 499.790 488.590 500.000 ;
        RECT 488.390 499.470 488.650 499.790 ;
        RECT 489.540 497.605 489.800 497.750 ;
        RECT 489.530 497.235 489.810 497.605 ;
        RECT 489.600 474.290 489.740 497.235 ;
        RECT 483.100 473.970 483.360 474.290 ;
        RECT 489.540 473.970 489.800 474.290 ;
        RECT 483.160 40.450 483.300 473.970 ;
        RECT 483.100 40.130 483.360 40.450 ;
        RECT 1026.360 40.130 1026.620 40.450 ;
        RECT 1026.420 2.400 1026.560 40.130 ;
        RECT 1026.210 -4.800 1026.770 2.400 ;
      LAYER via2 ;
        RECT 534.150 759.760 534.430 760.040 ;
        RECT 489.530 497.280 489.810 497.560 ;
      LAYER met3 ;
        RECT 418.870 760.050 419.250 760.060 ;
        RECT 534.125 760.050 534.455 760.065 ;
        RECT 418.870 759.750 534.455 760.050 ;
        RECT 418.870 759.740 419.250 759.750 ;
        RECT 534.125 759.735 534.455 759.750 ;
        RECT 418.870 500.290 419.250 500.300 ;
        RECT 418.870 499.990 444.050 500.290 ;
        RECT 418.870 499.980 419.250 499.990 ;
        RECT 443.750 497.570 444.050 499.990 ;
        RECT 489.505 497.570 489.835 497.585 ;
        RECT 443.750 497.270 489.835 497.570 ;
        RECT 489.505 497.255 489.835 497.270 ;
      LAYER via3 ;
        RECT 418.900 759.740 419.220 760.060 ;
        RECT 418.900 499.980 419.220 500.300 ;
      LAYER met4 ;
        RECT 418.895 759.735 419.225 760.065 ;
        RECT 418.910 500.305 419.210 759.735 ;
        RECT 418.895 499.975 419.225 500.305 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.570 761.160 540.890 761.220 ;
        RECT 540.570 761.020 590.020 761.160 ;
        RECT 540.570 760.960 540.890 761.020 ;
        RECT 589.880 760.820 590.020 761.020 ;
        RECT 642.230 760.820 642.550 760.880 ;
        RECT 589.880 760.680 642.550 760.820 ;
        RECT 642.230 760.620 642.550 760.680 ;
        RECT 489.740 499.500 490.060 499.760 ;
        RECT 489.830 498.060 489.970 499.500 ;
        RECT 489.830 497.860 490.290 498.060 ;
        RECT 489.970 497.800 490.290 497.860 ;
        RECT 489.510 471.480 489.830 471.540 ;
        RECT 492.270 471.480 492.590 471.540 ;
        RECT 489.510 471.340 492.590 471.480 ;
        RECT 489.510 471.280 489.830 471.340 ;
        RECT 492.270 471.280 492.590 471.340 ;
        RECT 492.270 441.560 492.590 441.620 ;
        RECT 642.230 441.560 642.550 441.620 ;
        RECT 1041.970 441.560 1042.290 441.620 ;
        RECT 492.270 441.420 1042.290 441.560 ;
        RECT 492.270 441.360 492.590 441.420 ;
        RECT 642.230 441.360 642.550 441.420 ;
        RECT 1041.970 441.360 1042.290 441.420 ;
      LAYER via ;
        RECT 540.600 760.960 540.860 761.220 ;
        RECT 642.260 760.620 642.520 760.880 ;
        RECT 489.770 499.500 490.030 499.760 ;
        RECT 490.000 497.800 490.260 498.060 ;
        RECT 489.540 471.280 489.800 471.540 ;
        RECT 492.300 471.280 492.560 471.540 ;
        RECT 492.300 441.360 492.560 441.620 ;
        RECT 642.260 441.360 642.520 441.620 ;
        RECT 1042.000 441.360 1042.260 441.620 ;
      LAYER met2 ;
        RECT 540.600 760.930 540.860 761.250 ;
        RECT 540.660 750.000 540.800 760.930 ;
        RECT 642.260 760.590 642.520 760.910 ;
        RECT 540.390 749.630 540.800 750.000 ;
        RECT 540.390 746.000 540.670 749.630 ;
        RECT 489.790 500.000 490.070 504.000 ;
        RECT 489.830 499.790 489.970 500.000 ;
        RECT 489.770 499.470 490.030 499.790 ;
        RECT 490.000 497.770 490.260 498.090 ;
        RECT 490.060 473.690 490.200 497.770 ;
        RECT 489.600 473.550 490.200 473.690 ;
        RECT 489.600 471.570 489.740 473.550 ;
        RECT 489.540 471.250 489.800 471.570 ;
        RECT 492.300 471.250 492.560 471.570 ;
        RECT 492.360 441.650 492.500 471.250 ;
        RECT 642.320 441.650 642.460 760.590 ;
        RECT 492.300 441.330 492.560 441.650 ;
        RECT 642.260 441.330 642.520 441.650 ;
        RECT 1042.000 441.330 1042.260 441.650 ;
        RECT 1042.060 17.410 1042.200 441.330 ;
        RECT 1042.060 17.270 1043.120 17.410 ;
        RECT 1042.980 2.400 1043.120 17.270 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.550 764.560 546.870 764.620 ;
        RECT 643.610 764.560 643.930 764.620 ;
        RECT 546.550 764.420 643.930 764.560 ;
        RECT 546.550 764.360 546.870 764.420 ;
        RECT 643.610 764.360 643.930 764.420 ;
        RECT 491.120 499.500 491.440 499.760 ;
        RECT 491.210 498.340 491.350 499.500 ;
        RECT 492.270 498.340 492.590 498.400 ;
        RECT 491.210 498.200 492.590 498.340 ;
        RECT 492.270 498.140 492.590 498.200 ;
        RECT 492.270 489.160 492.590 489.220 ;
        RECT 494.110 489.160 494.430 489.220 ;
        RECT 492.270 489.020 494.430 489.160 ;
        RECT 492.270 488.960 492.590 489.020 ;
        RECT 494.110 488.960 494.430 489.020 ;
        RECT 494.110 455.160 494.430 455.220 ;
        RECT 643.610 455.160 643.930 455.220 ;
        RECT 494.110 455.020 643.930 455.160 ;
        RECT 494.110 454.960 494.430 455.020 ;
        RECT 643.610 454.960 643.930 455.020 ;
        RECT 643.610 453.120 643.930 453.180 ;
        RECT 1055.770 453.120 1056.090 453.180 ;
        RECT 643.610 452.980 1056.090 453.120 ;
        RECT 643.610 452.920 643.930 452.980 ;
        RECT 1055.770 452.920 1056.090 452.980 ;
      LAYER via ;
        RECT 546.580 764.360 546.840 764.620 ;
        RECT 643.640 764.360 643.900 764.620 ;
        RECT 491.150 499.500 491.410 499.760 ;
        RECT 492.300 498.140 492.560 498.400 ;
        RECT 492.300 488.960 492.560 489.220 ;
        RECT 494.140 488.960 494.400 489.220 ;
        RECT 494.140 454.960 494.400 455.220 ;
        RECT 643.640 454.960 643.900 455.220 ;
        RECT 643.640 452.920 643.900 453.180 ;
        RECT 1055.800 452.920 1056.060 453.180 ;
      LAYER met2 ;
        RECT 546.580 764.330 546.840 764.650 ;
        RECT 643.640 764.330 643.900 764.650 ;
        RECT 545.910 749.770 546.190 750.000 ;
        RECT 546.640 749.770 546.780 764.330 ;
        RECT 545.910 749.630 546.780 749.770 ;
        RECT 545.910 746.000 546.190 749.630 ;
        RECT 491.170 500.000 491.450 504.000 ;
        RECT 491.210 499.790 491.350 500.000 ;
        RECT 491.150 499.470 491.410 499.790 ;
        RECT 492.300 498.110 492.560 498.430 ;
        RECT 492.360 489.250 492.500 498.110 ;
        RECT 492.300 488.930 492.560 489.250 ;
        RECT 494.140 488.930 494.400 489.250 ;
        RECT 494.200 455.250 494.340 488.930 ;
        RECT 643.700 455.250 643.840 764.330 ;
        RECT 494.140 454.930 494.400 455.250 ;
        RECT 643.640 454.930 643.900 455.250 ;
        RECT 643.700 453.210 643.840 454.930 ;
        RECT 643.640 452.890 643.900 453.210 ;
        RECT 1055.800 452.890 1056.060 453.210 ;
        RECT 1055.860 82.870 1056.000 452.890 ;
        RECT 1055.860 82.730 1059.680 82.870 ;
        RECT 1059.540 2.400 1059.680 82.730 ;
        RECT 1059.330 -4.800 1059.890 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 494.110 40.020 494.430 40.080 ;
        RECT 1076.010 40.020 1076.330 40.080 ;
        RECT 494.110 39.880 1076.330 40.020 ;
        RECT 494.110 39.820 494.430 39.880 ;
        RECT 1076.010 39.820 1076.330 39.880 ;
      LAYER via ;
        RECT 494.140 39.820 494.400 40.080 ;
        RECT 1076.040 39.820 1076.300 40.080 ;
      LAYER met2 ;
        RECT 551.630 763.115 551.910 763.485 ;
        RECT 551.700 750.000 551.840 763.115 ;
        RECT 551.430 749.630 551.840 750.000 ;
        RECT 551.430 746.000 551.710 749.630 ;
        RECT 492.550 500.000 492.830 504.000 ;
        RECT 492.590 499.815 492.730 500.000 ;
        RECT 492.520 499.445 492.800 499.815 ;
        RECT 493.210 497.915 493.490 498.285 ;
        RECT 493.280 488.765 493.420 497.915 ;
        RECT 493.210 488.395 493.490 488.765 ;
        RECT 493.280 448.570 493.420 488.395 ;
        RECT 493.280 448.430 494.800 448.570 ;
        RECT 494.660 420.970 494.800 448.430 ;
        RECT 494.200 420.830 494.800 420.970 ;
        RECT 494.200 40.110 494.340 420.830 ;
        RECT 494.140 39.790 494.400 40.110 ;
        RECT 1076.040 39.790 1076.300 40.110 ;
        RECT 1076.100 2.400 1076.240 39.790 ;
        RECT 1075.890 -4.800 1076.450 2.400 ;
      LAYER via2 ;
        RECT 551.630 763.160 551.910 763.440 ;
        RECT 492.520 499.490 492.800 499.770 ;
        RECT 493.210 497.960 493.490 498.240 ;
        RECT 493.210 488.440 493.490 488.720 ;
      LAYER met3 ;
        RECT 551.605 763.450 551.935 763.465 ;
        RECT 612.990 763.450 613.370 763.460 ;
        RECT 551.605 763.150 613.370 763.450 ;
        RECT 551.605 763.135 551.935 763.150 ;
        RECT 612.990 763.140 613.370 763.150 ;
        RECT 492.495 499.465 492.825 499.795 ;
        RECT 492.510 498.250 492.810 499.465 ;
        RECT 493.185 498.250 493.515 498.265 ;
        RECT 492.510 497.950 493.515 498.250 ;
        RECT 493.185 497.935 493.515 497.950 ;
        RECT 493.185 488.730 493.515 488.745 ;
        RECT 614.830 488.730 615.210 488.740 ;
        RECT 493.185 488.430 615.210 488.730 ;
        RECT 493.185 488.415 493.515 488.430 ;
        RECT 614.830 488.420 615.210 488.430 ;
      LAYER via3 ;
        RECT 613.020 763.140 613.340 763.460 ;
        RECT 614.860 488.420 615.180 488.740 ;
      LAYER met4 ;
        RECT 613.015 763.135 613.345 763.465 ;
        RECT 613.030 545.250 613.330 763.135 ;
        RECT 613.030 544.950 615.170 545.250 ;
        RECT 614.870 488.745 615.170 544.950 ;
        RECT 614.855 488.415 615.185 488.745 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 557.130 760.820 557.450 760.880 ;
        RECT 588.870 760.820 589.190 760.880 ;
        RECT 557.130 760.680 589.190 760.820 ;
        RECT 557.130 760.620 557.450 760.680 ;
        RECT 588.870 760.620 589.190 760.680 ;
        RECT 588.870 759.460 589.190 759.520 ;
        RECT 643.150 759.460 643.470 759.520 ;
        RECT 588.870 759.320 643.470 759.460 ;
        RECT 588.870 759.260 589.190 759.320 ;
        RECT 643.150 759.260 643.470 759.320 ;
        RECT 492.730 487.800 493.050 487.860 ;
        RECT 495.950 487.800 496.270 487.860 ;
        RECT 492.730 487.660 496.270 487.800 ;
        RECT 492.730 487.600 493.050 487.660 ;
        RECT 495.950 487.600 496.270 487.660 ;
        RECT 492.730 448.360 493.050 448.420 ;
        RECT 641.770 448.360 642.090 448.420 ;
        RECT 492.730 448.220 642.090 448.360 ;
        RECT 492.730 448.160 493.050 448.220 ;
        RECT 641.770 448.160 642.090 448.220 ;
        RECT 641.770 447.000 642.090 447.060 ;
        RECT 643.150 447.000 643.470 447.060 ;
        RECT 1090.270 447.000 1090.590 447.060 ;
        RECT 641.770 446.860 1090.590 447.000 ;
        RECT 641.770 446.800 642.090 446.860 ;
        RECT 643.150 446.800 643.470 446.860 ;
        RECT 1090.270 446.800 1090.590 446.860 ;
      LAYER via ;
        RECT 557.160 760.620 557.420 760.880 ;
        RECT 588.900 760.620 589.160 760.880 ;
        RECT 588.900 759.260 589.160 759.520 ;
        RECT 643.180 759.260 643.440 759.520 ;
        RECT 492.760 487.600 493.020 487.860 ;
        RECT 495.980 487.600 496.240 487.860 ;
        RECT 492.760 448.160 493.020 448.420 ;
        RECT 641.800 448.160 642.060 448.420 ;
        RECT 641.800 446.800 642.060 447.060 ;
        RECT 643.180 446.800 643.440 447.060 ;
        RECT 1090.300 446.800 1090.560 447.060 ;
      LAYER met2 ;
        RECT 557.160 760.590 557.420 760.910 ;
        RECT 588.900 760.590 589.160 760.910 ;
        RECT 557.220 750.000 557.360 760.590 ;
        RECT 588.960 759.550 589.100 760.590 ;
        RECT 588.900 759.230 589.160 759.550 ;
        RECT 643.180 759.230 643.440 759.550 ;
        RECT 556.950 749.630 557.360 750.000 ;
        RECT 556.950 746.000 557.230 749.630 ;
        RECT 493.930 500.000 494.210 504.000 ;
        RECT 493.970 499.645 494.110 500.000 ;
        RECT 493.900 499.275 494.180 499.645 ;
        RECT 495.970 498.595 496.250 498.965 ;
        RECT 496.040 487.890 496.180 498.595 ;
        RECT 492.760 487.570 493.020 487.890 ;
        RECT 495.980 487.570 496.240 487.890 ;
        RECT 492.820 448.450 492.960 487.570 ;
        RECT 492.760 448.130 493.020 448.450 ;
        RECT 641.800 448.130 642.060 448.450 ;
        RECT 641.860 447.090 642.000 448.130 ;
        RECT 643.240 447.090 643.380 759.230 ;
        RECT 641.800 446.770 642.060 447.090 ;
        RECT 643.180 446.770 643.440 447.090 ;
        RECT 1090.300 446.770 1090.560 447.090 ;
        RECT 1090.360 82.870 1090.500 446.770 ;
        RECT 1090.360 82.730 1092.800 82.870 ;
        RECT 1092.660 2.400 1092.800 82.730 ;
        RECT 1092.450 -4.800 1093.010 2.400 ;
      LAYER via2 ;
        RECT 493.900 499.320 494.180 499.600 ;
        RECT 495.970 498.640 496.250 498.920 ;
      LAYER met3 ;
        RECT 493.875 499.610 494.205 499.625 ;
        RECT 493.875 499.310 496.260 499.610 ;
        RECT 493.875 499.295 494.205 499.310 ;
        RECT 495.960 498.945 496.260 499.310 ;
        RECT 495.945 498.615 496.275 498.945 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 495.120 499.900 498.480 500.040 ;
        RECT 495.120 499.420 495.260 499.900 ;
        RECT 495.030 499.160 495.350 499.420 ;
        RECT 498.340 499.080 498.480 499.900 ;
        RECT 498.250 498.820 498.570 499.080 ;
        RECT 490.430 473.520 490.750 473.580 ;
        RECT 496.410 473.520 496.730 473.580 ;
        RECT 490.430 473.380 496.730 473.520 ;
        RECT 490.430 473.320 490.750 473.380 ;
        RECT 496.410 473.320 496.730 473.380 ;
        RECT 496.410 39.680 496.730 39.740 ;
        RECT 1109.130 39.680 1109.450 39.740 ;
        RECT 496.410 39.540 1109.450 39.680 ;
        RECT 496.410 39.480 496.730 39.540 ;
        RECT 1109.130 39.480 1109.450 39.540 ;
      LAYER via ;
        RECT 495.060 499.160 495.320 499.420 ;
        RECT 498.280 498.820 498.540 499.080 ;
        RECT 490.460 473.320 490.720 473.580 ;
        RECT 496.440 473.320 496.700 473.580 ;
        RECT 496.440 39.480 496.700 39.740 ;
        RECT 1109.160 39.480 1109.420 39.740 ;
      LAYER met2 ;
        RECT 563.130 759.715 563.410 760.085 ;
        RECT 562.470 749.770 562.750 750.000 ;
        RECT 563.200 749.770 563.340 759.715 ;
        RECT 562.470 749.630 563.340 749.770 ;
        RECT 562.470 746.000 562.750 749.630 ;
        RECT 495.310 500.000 495.590 504.000 ;
        RECT 495.350 499.530 495.490 500.000 ;
        RECT 495.120 499.450 495.490 499.530 ;
        RECT 495.060 499.390 495.490 499.450 ;
        RECT 495.060 499.130 495.320 499.390 ;
        RECT 498.280 498.965 498.540 499.110 ;
        RECT 498.270 498.595 498.550 498.965 ;
        RECT 490.450 484.995 490.730 485.365 ;
        RECT 490.520 473.610 490.660 484.995 ;
        RECT 490.460 473.290 490.720 473.610 ;
        RECT 496.440 473.290 496.700 473.610 ;
        RECT 496.500 39.770 496.640 473.290 ;
        RECT 496.440 39.450 496.700 39.770 ;
        RECT 1109.160 39.450 1109.420 39.770 ;
        RECT 1109.220 2.400 1109.360 39.450 ;
        RECT 1109.010 -4.800 1109.570 2.400 ;
      LAYER via2 ;
        RECT 563.130 759.760 563.410 760.040 ;
        RECT 498.270 498.640 498.550 498.920 ;
        RECT 490.450 485.040 490.730 485.320 ;
      LAYER met3 ;
        RECT 563.105 760.050 563.435 760.065 ;
        RECT 622.190 760.050 622.570 760.060 ;
        RECT 563.105 759.750 622.570 760.050 ;
        RECT 563.105 759.735 563.435 759.750 ;
        RECT 622.190 759.740 622.570 759.750 ;
        RECT 498.910 500.970 499.290 500.980 ;
        RECT 622.190 500.970 622.570 500.980 ;
        RECT 498.910 500.670 559.050 500.970 ;
        RECT 498.910 500.660 499.290 500.670 ;
        RECT 558.750 500.290 559.050 500.670 ;
        RECT 579.450 500.670 622.570 500.970 ;
        RECT 579.450 500.290 579.750 500.670 ;
        RECT 622.190 500.660 622.570 500.670 ;
        RECT 558.750 499.990 579.750 500.290 ;
        RECT 498.245 498.930 498.575 498.945 ;
        RECT 498.910 498.930 499.290 498.940 ;
        RECT 498.245 498.630 499.290 498.930 ;
        RECT 498.245 498.615 498.575 498.630 ;
        RECT 498.910 498.620 499.290 498.630 ;
        RECT 490.425 485.330 490.755 485.345 ;
        RECT 498.910 485.330 499.290 485.340 ;
        RECT 490.425 485.030 499.290 485.330 ;
        RECT 490.425 485.015 490.755 485.030 ;
        RECT 498.910 485.020 499.290 485.030 ;
      LAYER via3 ;
        RECT 622.220 759.740 622.540 760.060 ;
        RECT 498.940 500.660 499.260 500.980 ;
        RECT 622.220 500.660 622.540 500.980 ;
        RECT 498.940 498.620 499.260 498.940 ;
        RECT 498.940 485.020 499.260 485.340 ;
      LAYER met4 ;
        RECT 622.215 759.735 622.545 760.065 ;
        RECT 622.230 500.985 622.530 759.735 ;
        RECT 498.935 500.655 499.265 500.985 ;
        RECT 622.215 500.655 622.545 500.985 ;
        RECT 498.950 498.945 499.250 500.655 ;
        RECT 498.935 498.615 499.265 498.945 ;
        RECT 498.950 485.345 499.250 498.615 ;
        RECT 498.935 485.015 499.265 485.345 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.170 759.800 568.490 759.860 ;
        RECT 644.530 759.800 644.850 759.860 ;
        RECT 568.170 759.660 644.850 759.800 ;
        RECT 568.170 759.600 568.490 759.660 ;
        RECT 644.530 759.600 644.850 759.660 ;
        RECT 497.330 460.600 497.650 460.660 ;
        RECT 644.530 460.600 644.850 460.660 ;
        RECT 1124.770 460.600 1125.090 460.660 ;
        RECT 497.330 460.460 1125.090 460.600 ;
        RECT 497.330 460.400 497.650 460.460 ;
        RECT 644.530 460.400 644.850 460.460 ;
        RECT 1124.770 460.400 1125.090 460.460 ;
      LAYER via ;
        RECT 568.200 759.600 568.460 759.860 ;
        RECT 644.560 759.600 644.820 759.860 ;
        RECT 497.360 460.400 497.620 460.660 ;
        RECT 644.560 460.400 644.820 460.660 ;
        RECT 1124.800 460.400 1125.060 460.660 ;
      LAYER met2 ;
        RECT 568.200 759.570 568.460 759.890 ;
        RECT 644.560 759.570 644.820 759.890 ;
        RECT 568.260 750.000 568.400 759.570 ;
        RECT 567.990 749.630 568.400 750.000 ;
        RECT 567.990 746.000 568.270 749.630 ;
        RECT 496.690 500.000 496.970 504.000 ;
        RECT 496.730 498.680 496.870 500.000 ;
        RECT 496.730 498.540 497.560 498.680 ;
        RECT 497.420 460.690 497.560 498.540 ;
        RECT 644.620 460.690 644.760 759.570 ;
        RECT 497.360 460.370 497.620 460.690 ;
        RECT 644.560 460.370 644.820 460.690 ;
        RECT 1124.800 460.370 1125.060 460.690 ;
        RECT 1124.860 17.410 1125.000 460.370 ;
        RECT 1124.860 17.270 1125.920 17.410 ;
        RECT 1125.780 2.400 1125.920 17.270 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 762.520 574.470 762.580 ;
        RECT 590.250 762.520 590.570 762.580 ;
        RECT 574.150 762.380 590.570 762.520 ;
        RECT 574.150 762.320 574.470 762.380 ;
        RECT 590.250 762.320 590.570 762.380 ;
        RECT 590.250 761.160 590.570 761.220 ;
        RECT 642.690 761.160 643.010 761.220 ;
        RECT 590.250 761.020 643.010 761.160 ;
        RECT 590.250 760.960 590.570 761.020 ;
        RECT 642.690 760.960 643.010 761.020 ;
        RECT 498.020 500.380 498.340 500.440 ;
        RECT 498.020 500.240 499.170 500.380 ;
        RECT 498.020 500.180 498.340 500.240 ;
        RECT 499.030 498.000 499.170 500.240 ;
        RECT 499.630 498.000 499.950 498.060 ;
        RECT 499.030 497.860 499.950 498.000 ;
        RECT 499.630 497.800 499.950 497.860 ;
        RECT 499.630 441.220 499.950 441.280 ;
        RECT 642.690 441.220 643.010 441.280 ;
        RECT 1138.570 441.220 1138.890 441.280 ;
        RECT 499.630 441.080 1138.890 441.220 ;
        RECT 499.630 441.020 499.950 441.080 ;
        RECT 642.690 441.020 643.010 441.080 ;
        RECT 1138.570 441.020 1138.890 441.080 ;
      LAYER via ;
        RECT 574.180 762.320 574.440 762.580 ;
        RECT 590.280 762.320 590.540 762.580 ;
        RECT 590.280 760.960 590.540 761.220 ;
        RECT 642.720 760.960 642.980 761.220 ;
        RECT 498.050 500.180 498.310 500.440 ;
        RECT 499.660 497.800 499.920 498.060 ;
        RECT 499.660 441.020 499.920 441.280 ;
        RECT 642.720 441.020 642.980 441.280 ;
        RECT 1138.600 441.020 1138.860 441.280 ;
      LAYER met2 ;
        RECT 574.180 762.290 574.440 762.610 ;
        RECT 590.280 762.290 590.540 762.610 ;
        RECT 573.510 749.770 573.790 750.000 ;
        RECT 574.240 749.770 574.380 762.290 ;
        RECT 590.340 761.250 590.480 762.290 ;
        RECT 590.280 760.930 590.540 761.250 ;
        RECT 642.720 760.930 642.980 761.250 ;
        RECT 573.510 749.630 574.380 749.770 ;
        RECT 573.510 746.000 573.790 749.630 ;
        RECT 498.070 500.470 498.350 504.000 ;
        RECT 498.050 500.150 498.350 500.470 ;
        RECT 498.070 500.000 498.350 500.150 ;
        RECT 499.660 497.770 499.920 498.090 ;
        RECT 499.720 441.310 499.860 497.770 ;
        RECT 642.780 441.310 642.920 760.930 ;
        RECT 499.660 440.990 499.920 441.310 ;
        RECT 642.720 440.990 642.980 441.310 ;
        RECT 1138.600 440.990 1138.860 441.310 ;
        RECT 1138.660 82.870 1138.800 440.990 ;
        RECT 1138.660 82.730 1142.480 82.870 ;
        RECT 1142.340 2.400 1142.480 82.730 ;
        RECT 1142.130 -4.800 1142.690 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.210 761.500 579.530 761.560 ;
        RECT 639.930 761.500 640.250 761.560 ;
        RECT 579.210 761.360 640.250 761.500 ;
        RECT 579.210 761.300 579.530 761.360 ;
        RECT 639.930 761.300 640.250 761.360 ;
        RECT 545.030 502.960 552.070 503.100 ;
        RECT 545.030 501.060 545.170 502.960 ;
        RECT 551.930 502.760 552.070 502.960 ;
        RECT 551.930 502.620 579.670 502.760 ;
        RECT 501.790 500.920 545.170 501.060 ;
        RECT 579.530 501.060 579.670 502.620 ;
        RECT 593.330 501.260 600.370 501.400 ;
        RECT 593.330 501.060 593.470 501.260 ;
        RECT 579.530 500.920 593.470 501.060 ;
        RECT 600.230 501.060 600.370 501.260 ;
        RECT 600.230 500.920 627.970 501.060 ;
        RECT 500.090 497.320 500.410 497.380 ;
        RECT 501.790 497.320 501.930 500.920 ;
        RECT 627.830 500.720 627.970 500.920 ;
        RECT 639.930 500.720 640.250 500.780 ;
        RECT 627.830 500.580 640.250 500.720 ;
        RECT 639.930 500.520 640.250 500.580 ;
        RECT 500.090 497.180 501.930 497.320 ;
        RECT 500.090 497.120 500.410 497.180 ;
        RECT 500.090 472.840 500.410 472.900 ;
        RECT 503.310 472.840 503.630 472.900 ;
        RECT 500.090 472.700 503.630 472.840 ;
        RECT 500.090 472.640 500.410 472.700 ;
        RECT 503.310 472.640 503.630 472.700 ;
        RECT 503.310 39.000 503.630 39.060 ;
        RECT 1158.810 39.000 1159.130 39.060 ;
        RECT 503.310 38.860 1159.130 39.000 ;
        RECT 503.310 38.800 503.630 38.860 ;
        RECT 1158.810 38.800 1159.130 38.860 ;
      LAYER via ;
        RECT 579.240 761.300 579.500 761.560 ;
        RECT 639.960 761.300 640.220 761.560 ;
        RECT 500.120 497.120 500.380 497.380 ;
        RECT 639.960 500.520 640.220 500.780 ;
        RECT 500.120 472.640 500.380 472.900 ;
        RECT 503.340 472.640 503.600 472.900 ;
        RECT 503.340 38.800 503.600 39.060 ;
        RECT 1158.840 38.800 1159.100 39.060 ;
      LAYER met2 ;
        RECT 579.240 761.270 579.500 761.590 ;
        RECT 639.960 761.270 640.220 761.590 ;
        RECT 579.300 750.000 579.440 761.270 ;
        RECT 579.030 749.630 579.440 750.000 ;
        RECT 579.030 746.000 579.310 749.630 ;
        RECT 499.450 500.000 499.730 504.000 ;
        RECT 640.020 500.810 640.160 761.270 ;
        RECT 639.960 500.490 640.220 500.810 ;
        RECT 499.490 498.850 499.630 500.000 ;
        RECT 499.490 498.710 500.320 498.850 ;
        RECT 500.180 497.410 500.320 498.710 ;
        RECT 500.120 497.090 500.380 497.410 ;
        RECT 500.180 472.930 500.320 497.090 ;
        RECT 500.120 472.610 500.380 472.930 ;
        RECT 503.340 472.610 503.600 472.930 ;
        RECT 503.400 39.090 503.540 472.610 ;
        RECT 503.340 38.770 503.600 39.090 ;
        RECT 1158.840 38.770 1159.100 39.090 ;
        RECT 1158.900 2.400 1159.040 38.770 ;
        RECT 1158.690 -4.800 1159.250 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.730 759.120 585.050 759.180 ;
        RECT 640.850 759.120 641.170 759.180 ;
        RECT 584.730 758.980 596.000 759.120 ;
        RECT 584.730 758.920 585.050 758.980 ;
        RECT 595.860 758.780 596.000 758.980 ;
        RECT 603.680 758.980 641.170 759.120 ;
        RECT 603.680 758.780 603.820 758.980 ;
        RECT 640.850 758.920 641.170 758.980 ;
        RECT 595.860 758.640 603.820 758.780 ;
        RECT 565.730 503.980 572.770 504.120 ;
        RECT 565.730 503.440 565.870 503.980 ;
        RECT 572.630 503.780 572.770 503.980 ;
        RECT 572.630 503.640 579.670 503.780 ;
        RECT 516.050 503.300 565.870 503.440 ;
        RECT 516.050 502.420 516.190 503.300 ;
        RECT 579.530 503.100 579.670 503.640 ;
        RECT 579.530 502.960 600.370 503.100 ;
        RECT 500.640 502.280 516.190 502.420 ;
        RECT 600.230 502.420 600.370 502.960 ;
        RECT 600.230 502.280 614.170 502.420 ;
        RECT 500.640 500.720 500.780 502.280 ;
        RECT 614.030 501.740 614.170 502.280 ;
        RECT 640.850 501.740 641.170 501.800 ;
        RECT 614.030 501.600 641.170 501.740 ;
        RECT 640.850 501.540 641.170 501.600 ;
        RECT 499.950 500.580 500.780 500.720 ;
        RECT 499.950 499.700 500.090 500.580 ;
        RECT 500.780 499.700 501.100 499.760 ;
        RECT 499.950 499.560 501.100 499.700 ;
        RECT 500.780 499.500 501.100 499.560 ;
        RECT 501.470 411.640 501.790 411.700 ;
        RECT 502.850 411.640 503.170 411.700 ;
        RECT 501.470 411.500 503.170 411.640 ;
        RECT 501.470 411.440 501.790 411.500 ;
        RECT 502.850 411.440 503.170 411.500 ;
        RECT 502.850 46.480 503.170 46.540 ;
        RECT 1175.370 46.480 1175.690 46.540 ;
        RECT 502.850 46.340 1175.690 46.480 ;
        RECT 502.850 46.280 503.170 46.340 ;
        RECT 1175.370 46.280 1175.690 46.340 ;
      LAYER via ;
        RECT 584.760 758.920 585.020 759.180 ;
        RECT 640.880 758.920 641.140 759.180 ;
        RECT 640.880 501.540 641.140 501.800 ;
        RECT 500.810 499.500 501.070 499.760 ;
        RECT 501.500 411.440 501.760 411.700 ;
        RECT 502.880 411.440 503.140 411.700 ;
        RECT 502.880 46.280 503.140 46.540 ;
        RECT 1175.400 46.280 1175.660 46.540 ;
      LAYER met2 ;
        RECT 584.760 758.890 585.020 759.210 ;
        RECT 640.880 758.890 641.140 759.210 ;
        RECT 584.820 750.000 584.960 758.890 ;
        RECT 584.550 749.630 584.960 750.000 ;
        RECT 584.550 746.000 584.830 749.630 ;
        RECT 500.830 500.000 501.110 504.000 ;
        RECT 640.940 501.830 641.080 758.890 ;
        RECT 640.880 501.510 641.140 501.830 ;
        RECT 500.870 499.790 501.010 500.000 ;
        RECT 500.810 499.470 501.070 499.790 ;
        RECT 500.870 499.020 501.010 499.470 ;
        RECT 500.870 498.880 502.160 499.020 ;
        RECT 502.020 483.070 502.160 498.880 ;
        RECT 501.560 482.930 502.160 483.070 ;
        RECT 501.560 411.730 501.700 482.930 ;
        RECT 501.500 411.410 501.760 411.730 ;
        RECT 502.880 411.410 503.140 411.730 ;
        RECT 502.940 46.570 503.080 411.410 ;
        RECT 502.880 46.250 503.140 46.570 ;
        RECT 1175.400 46.250 1175.660 46.570 ;
        RECT 1175.460 2.400 1175.600 46.250 ;
        RECT 1175.250 -4.800 1175.810 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 409.010 747.900 409.330 747.960 ;
        RECT 434.770 747.900 435.090 747.960 ;
        RECT 409.010 747.760 435.090 747.900 ;
        RECT 409.010 747.700 409.330 747.760 ;
        RECT 434.770 747.700 435.090 747.760 ;
        RECT 455.100 499.900 463.750 500.040 ;
        RECT 455.100 498.060 455.240 499.900 ;
        RECT 463.610 499.760 463.750 499.900 ;
        RECT 463.520 499.500 463.840 499.760 ;
        RECT 455.010 497.800 455.330 498.060 ;
        RECT 407.630 486.100 407.950 486.160 ;
        RECT 455.010 486.100 455.330 486.160 ;
        RECT 468.350 486.100 468.670 486.160 ;
        RECT 407.630 485.960 468.670 486.100 ;
        RECT 407.630 485.900 407.950 485.960 ;
        RECT 455.010 485.900 455.330 485.960 ;
        RECT 468.350 485.900 468.670 485.960 ;
        RECT 462.830 471.140 463.150 471.200 ;
        RECT 468.350 471.140 468.670 471.200 ;
        RECT 462.830 471.000 468.670 471.140 ;
        RECT 462.830 470.940 463.150 471.000 ;
        RECT 468.350 470.940 468.670 471.000 ;
        RECT 462.830 448.020 463.150 448.080 ;
        RECT 724.570 448.020 724.890 448.080 ;
        RECT 462.830 447.880 724.890 448.020 ;
        RECT 462.830 447.820 463.150 447.880 ;
        RECT 724.570 447.820 724.890 447.880 ;
      LAYER via ;
        RECT 409.040 747.700 409.300 747.960 ;
        RECT 434.800 747.700 435.060 747.960 ;
        RECT 463.550 499.500 463.810 499.760 ;
        RECT 455.040 497.800 455.300 498.060 ;
        RECT 407.660 485.900 407.920 486.160 ;
        RECT 455.040 485.900 455.300 486.160 ;
        RECT 468.380 485.900 468.640 486.160 ;
        RECT 462.860 470.940 463.120 471.200 ;
        RECT 468.380 470.940 468.640 471.200 ;
        RECT 462.860 447.820 463.120 448.080 ;
        RECT 724.600 447.820 724.860 448.080 ;
      LAYER met2 ;
        RECT 409.040 747.670 409.300 747.990 ;
        RECT 434.800 747.730 435.060 747.990 ;
        RECT 435.510 747.730 435.790 750.000 ;
        RECT 434.800 747.670 435.790 747.730 ;
        RECT 409.100 522.085 409.240 747.670 ;
        RECT 434.860 747.590 435.790 747.670 ;
        RECT 435.510 746.000 435.790 747.590 ;
        RECT 407.650 521.715 407.930 522.085 ;
        RECT 409.030 521.715 409.310 522.085 ;
        RECT 407.720 486.190 407.860 521.715 ;
        RECT 463.570 500.000 463.850 504.000 ;
        RECT 463.610 499.790 463.750 500.000 ;
        RECT 463.550 499.470 463.810 499.790 ;
        RECT 455.040 497.770 455.300 498.090 ;
        RECT 455.100 486.190 455.240 497.770 ;
        RECT 407.660 485.870 407.920 486.190 ;
        RECT 455.040 485.870 455.300 486.190 ;
        RECT 468.380 485.870 468.640 486.190 ;
        RECT 468.440 471.230 468.580 485.870 ;
        RECT 462.860 470.910 463.120 471.230 ;
        RECT 468.380 470.910 468.640 471.230 ;
        RECT 462.920 448.110 463.060 470.910 ;
        RECT 462.860 447.790 463.120 448.110 ;
        RECT 724.600 447.790 724.860 448.110 ;
        RECT 724.660 82.870 724.800 447.790 ;
        RECT 724.660 82.730 728.480 82.870 ;
        RECT 728.340 2.400 728.480 82.730 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 407.650 521.760 407.930 522.040 ;
        RECT 409.030 521.760 409.310 522.040 ;
      LAYER met3 ;
        RECT 407.625 522.050 407.955 522.065 ;
        RECT 409.005 522.050 409.335 522.065 ;
        RECT 407.625 521.750 409.335 522.050 ;
        RECT 407.625 521.735 407.955 521.750 ;
        RECT 409.005 521.735 409.335 521.750 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.710 747.900 591.030 747.960 ;
        RECT 640.390 747.900 640.710 747.960 ;
        RECT 590.710 747.760 640.710 747.900 ;
        RECT 590.710 747.700 591.030 747.760 ;
        RECT 640.390 747.700 640.710 747.760 ;
        RECT 502.250 500.580 563.570 500.720 ;
        RECT 502.250 499.760 502.390 500.580 ;
        RECT 502.160 499.500 502.480 499.760 ;
        RECT 502.250 499.020 502.390 499.500 ;
        RECT 502.250 498.880 502.620 499.020 ;
        RECT 502.480 498.060 502.620 498.880 ;
        RECT 502.390 497.800 502.710 498.060 ;
        RECT 563.430 497.660 563.570 500.580 ;
        RECT 624.380 498.540 627.970 498.680 ;
        RECT 563.430 497.520 565.870 497.660 ;
        RECT 565.730 496.300 565.870 497.520 ;
        RECT 624.380 496.980 624.520 498.540 ;
        RECT 574.240 496.840 624.520 496.980 ;
        RECT 574.240 496.300 574.380 496.840 ;
        RECT 627.830 496.640 627.970 498.540 ;
        RECT 640.390 496.640 640.710 496.700 ;
        RECT 627.830 496.500 640.710 496.640 ;
        RECT 640.390 496.440 640.710 496.500 ;
        RECT 565.730 496.160 574.380 496.300 ;
        RECT 502.390 198.800 502.710 198.860 ;
        RECT 1186.870 198.800 1187.190 198.860 ;
        RECT 502.390 198.660 1187.190 198.800 ;
        RECT 502.390 198.600 502.710 198.660 ;
        RECT 1186.870 198.600 1187.190 198.660 ;
      LAYER via ;
        RECT 590.740 747.700 591.000 747.960 ;
        RECT 640.420 747.700 640.680 747.960 ;
        RECT 502.190 499.500 502.450 499.760 ;
        RECT 502.420 497.800 502.680 498.060 ;
        RECT 640.420 496.440 640.680 496.700 ;
        RECT 502.420 198.600 502.680 198.860 ;
        RECT 1186.900 198.600 1187.160 198.860 ;
      LAYER met2 ;
        RECT 590.070 747.730 590.350 750.000 ;
        RECT 590.740 747.730 591.000 747.990 ;
        RECT 590.070 747.670 591.000 747.730 ;
        RECT 640.420 747.670 640.680 747.990 ;
        RECT 590.070 747.590 590.940 747.670 ;
        RECT 590.070 746.000 590.350 747.590 ;
        RECT 502.210 500.000 502.490 504.000 ;
        RECT 502.250 499.790 502.390 500.000 ;
        RECT 502.190 499.470 502.450 499.790 ;
        RECT 502.420 497.770 502.680 498.090 ;
        RECT 502.480 476.170 502.620 497.770 ;
        RECT 640.480 496.730 640.620 747.670 ;
        RECT 640.420 496.410 640.680 496.730 ;
        RECT 502.480 476.030 503.080 476.170 ;
        RECT 502.940 473.010 503.080 476.030 ;
        RECT 502.020 472.870 503.080 473.010 ;
        RECT 502.020 471.820 502.160 472.870 ;
        RECT 502.020 471.680 502.620 471.820 ;
        RECT 502.480 434.770 502.620 471.680 ;
        RECT 502.020 434.630 502.620 434.770 ;
        RECT 502.020 386.470 502.160 434.630 ;
        RECT 502.020 386.330 502.620 386.470 ;
        RECT 502.480 198.890 502.620 386.330 ;
        RECT 502.420 198.570 502.680 198.890 ;
        RECT 1186.900 198.570 1187.160 198.890 ;
        RECT 1186.960 82.870 1187.100 198.570 ;
        RECT 1186.960 82.730 1192.160 82.870 ;
        RECT 1192.020 2.400 1192.160 82.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.540 500.180 503.860 500.440 ;
        RECT 503.630 500.040 503.770 500.180 ;
        RECT 503.630 499.900 509.980 500.040 ;
        RECT 509.840 497.720 509.980 499.900 ;
        RECT 509.750 497.460 510.070 497.720 ;
        RECT 590.710 487.800 591.030 487.860 ;
        RECT 579.530 487.660 591.030 487.800 ;
        RECT 509.750 487.120 510.070 487.180 ;
        RECT 579.530 487.120 579.670 487.660 ;
        RECT 590.710 487.600 591.030 487.660 ;
        RECT 509.750 486.980 579.670 487.120 ;
        RECT 509.750 486.920 510.070 486.980 ;
        RECT 590.710 485.420 591.030 485.480 ;
        RECT 598.990 485.420 599.310 485.480 ;
        RECT 590.710 485.280 599.310 485.420 ;
        RECT 590.710 485.220 591.030 485.280 ;
        RECT 598.990 485.220 599.310 485.280 ;
        RECT 598.990 446.660 599.310 446.720 ;
        RECT 649.130 446.660 649.450 446.720 ;
        RECT 1207.570 446.660 1207.890 446.720 ;
        RECT 598.990 446.520 1207.890 446.660 ;
        RECT 598.990 446.460 599.310 446.520 ;
        RECT 649.130 446.460 649.450 446.520 ;
        RECT 1207.570 446.460 1207.890 446.520 ;
      LAYER via ;
        RECT 503.570 500.180 503.830 500.440 ;
        RECT 509.780 497.460 510.040 497.720 ;
        RECT 509.780 486.920 510.040 487.180 ;
        RECT 590.740 487.600 591.000 487.860 ;
        RECT 590.740 485.220 591.000 485.480 ;
        RECT 599.020 485.220 599.280 485.480 ;
        RECT 599.020 446.460 599.280 446.720 ;
        RECT 649.160 446.460 649.420 446.720 ;
        RECT 1207.600 446.460 1207.860 446.720 ;
      LAYER met2 ;
        RECT 595.790 759.035 596.070 759.405 ;
        RECT 649.150 759.035 649.430 759.405 ;
        RECT 595.860 750.000 596.000 759.035 ;
        RECT 595.590 749.630 596.000 750.000 ;
        RECT 595.590 746.000 595.870 749.630 ;
        RECT 503.590 500.470 503.870 504.000 ;
        RECT 503.570 500.150 503.870 500.470 ;
        RECT 503.590 500.000 503.870 500.150 ;
        RECT 509.780 497.430 510.040 497.750 ;
        RECT 509.840 487.210 509.980 497.430 ;
        RECT 590.740 487.570 591.000 487.890 ;
        RECT 509.780 486.890 510.040 487.210 ;
        RECT 590.800 485.510 590.940 487.570 ;
        RECT 590.740 485.190 591.000 485.510 ;
        RECT 599.020 485.190 599.280 485.510 ;
        RECT 599.080 446.750 599.220 485.190 ;
        RECT 649.220 446.750 649.360 759.035 ;
        RECT 599.020 446.430 599.280 446.750 ;
        RECT 649.160 446.430 649.420 446.750 ;
        RECT 1207.600 446.430 1207.860 446.750 ;
        RECT 1207.660 17.410 1207.800 446.430 ;
        RECT 1207.660 17.270 1208.720 17.410 ;
        RECT 1208.580 2.400 1208.720 17.270 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
      LAYER via2 ;
        RECT 595.790 759.080 596.070 759.360 ;
        RECT 649.150 759.080 649.430 759.360 ;
      LAYER met3 ;
        RECT 595.765 759.370 596.095 759.385 ;
        RECT 649.125 759.370 649.455 759.385 ;
        RECT 595.765 759.070 649.455 759.370 ;
        RECT 595.765 759.055 596.095 759.070 ;
        RECT 649.125 759.055 649.455 759.070 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.990 433.060 507.310 433.120 ;
        RECT 1221.370 433.060 1221.690 433.120 ;
        RECT 506.990 432.920 1221.690 433.060 ;
        RECT 506.990 432.860 507.310 432.920 ;
        RECT 1221.370 432.860 1221.690 432.920 ;
      LAYER via ;
        RECT 507.020 432.860 507.280 433.120 ;
        RECT 1221.400 432.860 1221.660 433.120 ;
      LAYER met2 ;
        RECT 504.970 500.000 505.250 504.000 ;
        RECT 505.010 499.815 505.150 500.000 ;
        RECT 504.940 499.445 505.220 499.815 ;
        RECT 507.010 497.235 507.290 497.605 ;
        RECT 507.080 433.150 507.220 497.235 ;
        RECT 507.020 432.830 507.280 433.150 ;
        RECT 1221.400 432.830 1221.660 433.150 ;
        RECT 1221.460 82.870 1221.600 432.830 ;
        RECT 1221.460 82.730 1225.280 82.870 ;
        RECT 1225.140 2.400 1225.280 82.730 ;
        RECT 1224.930 -4.800 1225.490 2.400 ;
      LAYER via2 ;
        RECT 504.940 499.490 505.220 499.770 ;
        RECT 507.010 497.280 507.290 497.560 ;
      LAYER met3 ;
        RECT 504.915 499.780 505.245 499.795 ;
        RECT 504.915 499.465 505.460 499.780 ;
        RECT 505.160 497.570 505.460 499.465 ;
        RECT 506.985 497.570 507.315 497.585 ;
        RECT 505.160 497.270 507.315 497.570 ;
        RECT 506.985 497.255 507.315 497.270 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.300 499.500 506.620 499.760 ;
        RECT 506.390 498.060 506.530 499.500 ;
        RECT 506.390 497.860 506.850 498.060 ;
        RECT 506.530 497.800 506.850 497.860 ;
        RECT 506.530 432.720 506.850 432.780 ;
        RECT 1235.630 432.720 1235.950 432.780 ;
        RECT 506.530 432.580 1235.950 432.720 ;
        RECT 506.530 432.520 506.850 432.580 ;
        RECT 1235.630 432.520 1235.950 432.580 ;
        RECT 1235.630 19.620 1235.950 19.680 ;
        RECT 1241.610 19.620 1241.930 19.680 ;
        RECT 1235.630 19.480 1241.930 19.620 ;
        RECT 1235.630 19.420 1235.950 19.480 ;
        RECT 1241.610 19.420 1241.930 19.480 ;
      LAYER via ;
        RECT 506.330 499.500 506.590 499.760 ;
        RECT 506.560 497.800 506.820 498.060 ;
        RECT 506.560 432.520 506.820 432.780 ;
        RECT 1235.660 432.520 1235.920 432.780 ;
        RECT 1235.660 19.420 1235.920 19.680 ;
        RECT 1241.640 19.420 1241.900 19.680 ;
      LAYER met2 ;
        RECT 506.350 500.000 506.630 504.000 ;
        RECT 506.390 499.790 506.530 500.000 ;
        RECT 506.330 499.470 506.590 499.790 ;
        RECT 506.560 497.770 506.820 498.090 ;
        RECT 506.620 432.810 506.760 497.770 ;
        RECT 506.560 432.490 506.820 432.810 ;
        RECT 1235.660 432.490 1235.920 432.810 ;
        RECT 1235.720 19.710 1235.860 432.490 ;
        RECT 1235.660 19.390 1235.920 19.710 ;
        RECT 1241.640 19.390 1241.900 19.710 ;
        RECT 1241.700 2.400 1241.840 19.390 ;
        RECT 1241.490 -4.800 1242.050 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 507.680 499.020 508.000 499.080 ;
        RECT 507.680 498.880 508.600 499.020 ;
        RECT 507.680 498.820 508.000 498.880 ;
        RECT 507.450 498.000 507.770 498.060 ;
        RECT 508.460 498.000 508.600 498.880 ;
        RECT 507.450 497.860 508.600 498.000 ;
        RECT 507.450 497.800 507.770 497.860 ;
        RECT 507.450 440.880 507.770 440.940 ;
        RECT 1255.870 440.880 1256.190 440.940 ;
        RECT 507.450 440.740 1256.190 440.880 ;
        RECT 507.450 440.680 507.770 440.740 ;
        RECT 1255.870 440.680 1256.190 440.740 ;
      LAYER via ;
        RECT 507.710 498.820 507.970 499.080 ;
        RECT 507.480 497.800 507.740 498.060 ;
        RECT 507.480 440.680 507.740 440.940 ;
        RECT 1255.900 440.680 1256.160 440.940 ;
      LAYER met2 ;
        RECT 507.730 500.000 508.010 504.000 ;
        RECT 507.770 499.110 507.910 500.000 ;
        RECT 507.710 498.790 507.970 499.110 ;
        RECT 507.480 497.770 507.740 498.090 ;
        RECT 507.540 440.970 507.680 497.770 ;
        RECT 507.480 440.650 507.740 440.970 ;
        RECT 1255.900 440.650 1256.160 440.970 ;
        RECT 1255.960 82.870 1256.100 440.650 ;
        RECT 1255.960 82.730 1258.400 82.870 ;
        RECT 1258.260 2.400 1258.400 82.730 ;
        RECT 1258.050 -4.800 1258.610 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.110 500.000 509.390 504.000 ;
        RECT 509.150 499.815 509.290 500.000 ;
        RECT 509.080 499.445 509.360 499.815 ;
        RECT 508.850 491.115 509.130 491.485 ;
        RECT 508.920 478.565 509.060 491.115 ;
        RECT 508.850 478.195 509.130 478.565 ;
        RECT 1274.750 44.355 1275.030 44.725 ;
        RECT 1274.820 2.400 1274.960 44.355 ;
        RECT 1274.610 -4.800 1275.170 2.400 ;
      LAYER via2 ;
        RECT 509.080 499.490 509.360 499.770 ;
        RECT 508.850 491.160 509.130 491.440 ;
        RECT 508.850 478.240 509.130 478.520 ;
        RECT 1274.750 44.400 1275.030 44.680 ;
      LAYER met3 ;
        RECT 509.055 499.620 509.385 499.795 ;
        RECT 509.030 499.610 509.410 499.620 ;
        RECT 509.030 499.310 509.670 499.610 ;
        RECT 509.030 499.300 509.410 499.310 ;
        RECT 508.825 491.460 509.155 491.465 ;
        RECT 508.825 491.450 509.410 491.460 ;
        RECT 508.600 491.150 509.410 491.450 ;
        RECT 508.825 491.140 509.410 491.150 ;
        RECT 508.825 491.135 509.155 491.140 ;
        RECT 508.825 478.530 509.155 478.545 ;
        RECT 509.950 478.530 510.330 478.540 ;
        RECT 508.825 478.230 510.330 478.530 ;
        RECT 508.825 478.215 509.155 478.230 ;
        RECT 509.950 478.220 510.330 478.230 ;
        RECT 509.950 44.690 510.330 44.700 ;
        RECT 1274.725 44.690 1275.055 44.705 ;
        RECT 509.950 44.390 1275.055 44.690 ;
        RECT 509.950 44.380 510.330 44.390 ;
        RECT 1274.725 44.375 1275.055 44.390 ;
      LAYER via3 ;
        RECT 509.060 499.300 509.380 499.620 ;
        RECT 509.060 491.140 509.380 491.460 ;
        RECT 509.980 478.220 510.300 478.540 ;
        RECT 509.980 44.380 510.300 44.700 ;
      LAYER met4 ;
        RECT 509.055 499.295 509.385 499.625 ;
        RECT 509.070 491.465 509.370 499.295 ;
        RECT 509.055 491.135 509.385 491.465 ;
        RECT 509.975 478.215 510.305 478.545 ;
        RECT 509.990 44.705 510.290 478.215 ;
        RECT 509.975 44.375 510.305 44.705 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.440 499.700 510.760 499.760 ;
        RECT 510.300 499.500 510.760 499.700 ;
        RECT 510.300 499.080 510.440 499.500 ;
        RECT 510.210 498.820 510.530 499.080 ;
        RECT 510.210 491.880 510.530 491.940 ;
        RECT 516.190 491.880 516.510 491.940 ;
        RECT 510.210 491.740 516.510 491.880 ;
        RECT 510.210 491.680 510.530 491.740 ;
        RECT 516.190 491.680 516.510 491.740 ;
        RECT 516.190 446.320 516.510 446.380 ;
        RECT 1290.370 446.320 1290.690 446.380 ;
        RECT 516.190 446.180 1290.690 446.320 ;
        RECT 516.190 446.120 516.510 446.180 ;
        RECT 1290.370 446.120 1290.690 446.180 ;
      LAYER via ;
        RECT 510.470 499.500 510.730 499.760 ;
        RECT 510.240 498.820 510.500 499.080 ;
        RECT 510.240 491.680 510.500 491.940 ;
        RECT 516.220 491.680 516.480 491.940 ;
        RECT 516.220 446.120 516.480 446.380 ;
        RECT 1290.400 446.120 1290.660 446.380 ;
      LAYER met2 ;
        RECT 510.490 500.000 510.770 504.000 ;
        RECT 510.530 499.790 510.670 500.000 ;
        RECT 510.470 499.470 510.730 499.790 ;
        RECT 510.240 498.790 510.500 499.110 ;
        RECT 510.300 491.970 510.440 498.790 ;
        RECT 510.240 491.650 510.500 491.970 ;
        RECT 516.220 491.650 516.480 491.970 ;
        RECT 516.280 446.410 516.420 491.650 ;
        RECT 516.220 446.090 516.480 446.410 ;
        RECT 1290.400 446.090 1290.660 446.410 ;
        RECT 1290.460 17.410 1290.600 446.090 ;
        RECT 1290.460 17.270 1291.520 17.410 ;
        RECT 1291.380 2.400 1291.520 17.270 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.820 499.500 512.140 499.760 ;
        RECT 511.910 499.360 512.050 499.500 ;
        RECT 511.910 499.220 512.280 499.360 ;
        RECT 512.140 498.740 512.280 499.220 ;
        RECT 512.050 498.480 512.370 498.740 ;
        RECT 511.590 46.140 511.910 46.200 ;
        RECT 1307.850 46.140 1308.170 46.200 ;
        RECT 511.590 46.000 1308.170 46.140 ;
        RECT 511.590 45.940 511.910 46.000 ;
        RECT 1307.850 45.940 1308.170 46.000 ;
      LAYER via ;
        RECT 511.850 499.500 512.110 499.760 ;
        RECT 512.080 498.480 512.340 498.740 ;
        RECT 511.620 45.940 511.880 46.200 ;
        RECT 1307.880 45.940 1308.140 46.200 ;
      LAYER met2 ;
        RECT 511.870 500.000 512.150 504.000 ;
        RECT 511.910 499.790 512.050 500.000 ;
        RECT 511.850 499.470 512.110 499.790 ;
        RECT 512.080 498.450 512.340 498.770 ;
        RECT 512.140 455.470 512.280 498.450 ;
        RECT 511.680 455.330 512.280 455.470 ;
        RECT 511.680 46.230 511.820 455.330 ;
        RECT 511.620 45.910 511.880 46.230 ;
        RECT 1307.880 45.910 1308.140 46.230 ;
        RECT 1307.940 2.400 1308.080 45.910 ;
        RECT 1307.730 -4.800 1308.290 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 513.200 499.360 513.520 499.420 ;
        RECT 513.060 499.160 513.520 499.360 ;
        RECT 513.060 498.060 513.200 499.160 ;
        RECT 512.970 497.800 513.290 498.060 ;
        RECT 510.670 477.940 510.990 478.000 ;
        RECT 512.970 477.940 513.290 478.000 ;
        RECT 510.670 477.800 513.290 477.940 ;
        RECT 510.670 477.740 510.990 477.800 ;
        RECT 512.970 477.740 513.290 477.800 ;
        RECT 510.670 45.800 510.990 45.860 ;
        RECT 1324.410 45.800 1324.730 45.860 ;
        RECT 510.670 45.660 1324.730 45.800 ;
        RECT 510.670 45.600 510.990 45.660 ;
        RECT 1324.410 45.600 1324.730 45.660 ;
      LAYER via ;
        RECT 513.230 499.160 513.490 499.420 ;
        RECT 513.000 497.800 513.260 498.060 ;
        RECT 510.700 477.740 510.960 478.000 ;
        RECT 513.000 477.740 513.260 478.000 ;
        RECT 510.700 45.600 510.960 45.860 ;
        RECT 1324.440 45.600 1324.700 45.860 ;
      LAYER met2 ;
        RECT 513.250 500.000 513.530 504.000 ;
        RECT 513.290 499.450 513.430 500.000 ;
        RECT 513.230 499.130 513.490 499.450 ;
        RECT 513.000 497.770 513.260 498.090 ;
        RECT 513.060 478.030 513.200 497.770 ;
        RECT 510.700 477.710 510.960 478.030 ;
        RECT 513.000 477.710 513.260 478.030 ;
        RECT 510.760 45.890 510.900 477.710 ;
        RECT 510.700 45.570 510.960 45.890 ;
        RECT 1324.440 45.570 1324.700 45.890 ;
        RECT 1324.500 2.400 1324.640 45.570 ;
        RECT 1324.290 -4.800 1324.850 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 45.460 511.450 45.520 ;
        RECT 1340.970 45.460 1341.290 45.520 ;
        RECT 511.130 45.320 1341.290 45.460 ;
        RECT 511.130 45.260 511.450 45.320 ;
        RECT 1340.970 45.260 1341.290 45.320 ;
      LAYER via ;
        RECT 511.160 45.260 511.420 45.520 ;
        RECT 1341.000 45.260 1341.260 45.520 ;
      LAYER met2 ;
        RECT 514.630 500.000 514.910 504.000 ;
        RECT 514.670 499.020 514.810 500.000 ;
        RECT 514.440 498.965 514.810 499.020 ;
        RECT 514.370 498.880 514.810 498.965 ;
        RECT 514.370 498.595 514.650 498.880 ;
        RECT 511.610 497.235 511.890 497.605 ;
        RECT 511.680 476.410 511.820 497.235 ;
        RECT 511.220 476.270 511.820 476.410 ;
        RECT 511.220 45.550 511.360 476.270 ;
        RECT 511.160 45.230 511.420 45.550 ;
        RECT 1341.000 45.230 1341.260 45.550 ;
        RECT 1341.060 2.400 1341.200 45.230 ;
        RECT 1340.850 -4.800 1341.410 2.400 ;
      LAYER via2 ;
        RECT 514.370 498.640 514.650 498.920 ;
        RECT 511.610 497.280 511.890 497.560 ;
      LAYER met3 ;
        RECT 514.345 498.930 514.675 498.945 ;
        RECT 514.345 498.615 514.890 498.930 ;
        RECT 511.585 497.570 511.915 497.585 ;
        RECT 514.590 497.570 514.890 498.615 ;
        RECT 511.585 497.270 514.890 497.570 ;
        RECT 511.585 497.255 511.915 497.270 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.900 499.500 465.220 499.760 ;
        RECT 464.990 498.340 465.130 499.500 ;
        RECT 464.990 498.200 465.820 498.340 ;
        RECT 465.680 498.060 465.820 498.200 ;
        RECT 465.590 497.800 465.910 498.060 ;
        RECT 465.590 53.960 465.910 54.020 ;
        RECT 738.830 53.960 739.150 54.020 ;
        RECT 465.590 53.820 739.150 53.960 ;
        RECT 465.590 53.760 465.910 53.820 ;
        RECT 738.830 53.760 739.150 53.820 ;
        RECT 738.830 19.960 739.150 20.020 ;
        RECT 744.810 19.960 745.130 20.020 ;
        RECT 738.830 19.820 745.130 19.960 ;
        RECT 738.830 19.760 739.150 19.820 ;
        RECT 744.810 19.760 745.130 19.820 ;
      LAYER via ;
        RECT 464.930 499.500 465.190 499.760 ;
        RECT 465.620 497.800 465.880 498.060 ;
        RECT 465.620 53.760 465.880 54.020 ;
        RECT 738.860 53.760 739.120 54.020 ;
        RECT 738.860 19.760 739.120 20.020 ;
        RECT 744.840 19.760 745.100 20.020 ;
      LAYER met2 ;
        RECT 440.310 747.050 440.590 747.165 ;
        RECT 441.030 747.050 441.310 750.000 ;
        RECT 440.310 746.910 441.310 747.050 ;
        RECT 440.310 746.795 440.590 746.910 ;
        RECT 441.030 746.000 441.310 746.910 ;
        RECT 464.950 500.000 465.230 504.000 ;
        RECT 464.990 499.790 465.130 500.000 ;
        RECT 464.930 499.470 465.190 499.790 ;
        RECT 465.620 497.770 465.880 498.090 ;
        RECT 465.680 488.085 465.820 497.770 ;
        RECT 465.610 487.715 465.890 488.085 ;
        RECT 465.680 54.050 465.820 487.715 ;
        RECT 465.620 53.730 465.880 54.050 ;
        RECT 738.860 53.730 739.120 54.050 ;
        RECT 738.920 20.050 739.060 53.730 ;
        RECT 738.860 19.730 739.120 20.050 ;
        RECT 744.840 19.730 745.100 20.050 ;
        RECT 744.900 2.400 745.040 19.730 ;
        RECT 744.690 -4.800 745.250 2.400 ;
      LAYER via2 ;
        RECT 440.310 746.840 440.590 747.120 ;
        RECT 465.610 487.760 465.890 488.040 ;
      LAYER met3 ;
        RECT 419.790 747.130 420.170 747.140 ;
        RECT 440.285 747.130 440.615 747.145 ;
        RECT 419.790 746.830 440.615 747.130 ;
        RECT 419.790 746.820 420.170 746.830 ;
        RECT 440.285 746.815 440.615 746.830 ;
        RECT 419.790 488.050 420.170 488.060 ;
        RECT 465.585 488.050 465.915 488.065 ;
        RECT 419.790 487.750 465.915 488.050 ;
        RECT 419.790 487.740 420.170 487.750 ;
        RECT 465.585 487.735 465.915 487.750 ;
      LAYER via3 ;
        RECT 419.820 746.820 420.140 747.140 ;
        RECT 419.820 487.740 420.140 488.060 ;
      LAYER met4 ;
        RECT 419.815 746.815 420.145 747.145 ;
        RECT 419.830 488.065 420.130 746.815 ;
        RECT 419.815 487.735 420.145 488.065 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.010 500.000 516.290 504.000 ;
        RECT 516.050 498.340 516.190 500.000 ;
        RECT 516.050 498.200 516.420 498.340 ;
        RECT 516.280 492.560 516.420 498.200 ;
        RECT 515.820 492.420 516.420 492.560 ;
        RECT 515.820 458.845 515.960 492.420 ;
        RECT 515.750 458.475 516.030 458.845 ;
        RECT 1352.490 424.475 1352.770 424.845 ;
        RECT 1352.560 82.870 1352.700 424.475 ;
        RECT 1352.560 82.730 1357.760 82.870 ;
        RECT 1357.620 2.400 1357.760 82.730 ;
        RECT 1357.410 -4.800 1357.970 2.400 ;
      LAYER via2 ;
        RECT 515.750 458.520 516.030 458.800 ;
        RECT 1352.490 424.520 1352.770 424.800 ;
      LAYER met3 ;
        RECT 513.630 458.810 514.010 458.820 ;
        RECT 515.725 458.810 516.055 458.825 ;
        RECT 513.630 458.510 516.055 458.810 ;
        RECT 513.630 458.500 514.010 458.510 ;
        RECT 515.725 458.495 516.055 458.510 ;
        RECT 513.630 424.810 514.010 424.820 ;
        RECT 1352.465 424.810 1352.795 424.825 ;
        RECT 513.630 424.510 1352.795 424.810 ;
        RECT 513.630 424.500 514.010 424.510 ;
        RECT 1352.465 424.495 1352.795 424.510 ;
      LAYER via3 ;
        RECT 513.660 458.500 513.980 458.820 ;
        RECT 513.660 424.500 513.980 424.820 ;
      LAYER met4 ;
        RECT 513.655 458.495 513.985 458.825 ;
        RECT 513.670 424.825 513.970 458.495 ;
        RECT 513.655 424.495 513.985 424.825 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.340 499.500 517.660 499.760 ;
        RECT 517.430 498.060 517.570 499.500 ;
        RECT 517.110 497.860 517.570 498.060 ;
        RECT 517.110 497.800 517.430 497.860 ;
        RECT 517.110 464.000 517.430 464.060 ;
        RECT 521.250 464.000 521.570 464.060 ;
        RECT 517.110 463.860 521.570 464.000 ;
        RECT 517.110 463.800 517.430 463.860 ;
        RECT 521.250 463.800 521.570 463.860 ;
        RECT 521.250 432.380 521.570 432.440 ;
        RECT 1373.170 432.380 1373.490 432.440 ;
        RECT 521.250 432.240 1373.490 432.380 ;
        RECT 521.250 432.180 521.570 432.240 ;
        RECT 1373.170 432.180 1373.490 432.240 ;
      LAYER via ;
        RECT 517.370 499.500 517.630 499.760 ;
        RECT 517.140 497.800 517.400 498.060 ;
        RECT 517.140 463.800 517.400 464.060 ;
        RECT 521.280 463.800 521.540 464.060 ;
        RECT 521.280 432.180 521.540 432.440 ;
        RECT 1373.200 432.180 1373.460 432.440 ;
      LAYER met2 ;
        RECT 517.390 500.000 517.670 504.000 ;
        RECT 517.430 499.790 517.570 500.000 ;
        RECT 517.370 499.470 517.630 499.790 ;
        RECT 517.140 497.770 517.400 498.090 ;
        RECT 517.200 464.090 517.340 497.770 ;
        RECT 517.140 463.770 517.400 464.090 ;
        RECT 521.280 463.770 521.540 464.090 ;
        RECT 521.340 432.470 521.480 463.770 ;
        RECT 521.280 432.150 521.540 432.470 ;
        RECT 1373.200 432.150 1373.460 432.470 ;
        RECT 1373.260 17.410 1373.400 432.150 ;
        RECT 1373.260 17.270 1374.320 17.410 ;
        RECT 1374.180 2.400 1374.320 17.270 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.720 499.500 519.040 499.760 ;
        RECT 518.810 497.720 518.950 499.500 ;
        RECT 518.490 497.520 518.950 497.720 ;
        RECT 518.490 497.460 518.810 497.520 ;
        RECT 517.570 480.320 517.890 480.380 ;
        RECT 518.490 480.320 518.810 480.380 ;
        RECT 517.570 480.180 518.810 480.320 ;
        RECT 517.570 480.120 517.890 480.180 ;
        RECT 518.490 480.120 518.810 480.180 ;
        RECT 517.570 45.120 517.890 45.180 ;
        RECT 1390.650 45.120 1390.970 45.180 ;
        RECT 517.570 44.980 1390.970 45.120 ;
        RECT 517.570 44.920 517.890 44.980 ;
        RECT 1390.650 44.920 1390.970 44.980 ;
      LAYER via ;
        RECT 518.750 499.500 519.010 499.760 ;
        RECT 518.520 497.460 518.780 497.720 ;
        RECT 517.600 480.120 517.860 480.380 ;
        RECT 518.520 480.120 518.780 480.380 ;
        RECT 517.600 44.920 517.860 45.180 ;
        RECT 1390.680 44.920 1390.940 45.180 ;
      LAYER met2 ;
        RECT 518.770 500.000 519.050 504.000 ;
        RECT 518.810 499.790 518.950 500.000 ;
        RECT 518.750 499.470 519.010 499.790 ;
        RECT 518.520 497.430 518.780 497.750 ;
        RECT 518.580 480.410 518.720 497.430 ;
        RECT 517.600 480.090 517.860 480.410 ;
        RECT 518.520 480.090 518.780 480.410 ;
        RECT 517.660 45.210 517.800 480.090 ;
        RECT 517.600 44.890 517.860 45.210 ;
        RECT 1390.680 44.890 1390.940 45.210 ;
        RECT 1390.740 2.400 1390.880 44.890 ;
        RECT 1390.530 -4.800 1391.090 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.190 499.900 521.250 500.040 ;
        RECT 520.190 499.760 520.330 499.900 ;
        RECT 520.100 499.500 520.420 499.760 ;
        RECT 518.950 497.320 519.270 497.380 ;
        RECT 521.110 497.320 521.250 499.900 ;
        RECT 518.950 497.180 521.250 497.320 ;
        RECT 518.950 497.120 519.270 497.180 ;
        RECT 518.030 490.860 518.350 490.920 ;
        RECT 518.950 490.860 519.270 490.920 ;
        RECT 518.030 490.720 519.270 490.860 ;
        RECT 518.030 490.660 518.350 490.720 ;
        RECT 518.950 490.660 519.270 490.720 ;
        RECT 518.490 53.280 518.810 53.340 ;
        RECT 1401.230 53.280 1401.550 53.340 ;
        RECT 518.490 53.140 1401.550 53.280 ;
        RECT 518.490 53.080 518.810 53.140 ;
        RECT 1401.230 53.080 1401.550 53.140 ;
        RECT 1401.230 19.620 1401.550 19.680 ;
        RECT 1407.210 19.620 1407.530 19.680 ;
        RECT 1401.230 19.480 1407.530 19.620 ;
        RECT 1401.230 19.420 1401.550 19.480 ;
        RECT 1407.210 19.420 1407.530 19.480 ;
      LAYER via ;
        RECT 520.130 499.500 520.390 499.760 ;
        RECT 518.980 497.120 519.240 497.380 ;
        RECT 518.060 490.660 518.320 490.920 ;
        RECT 518.980 490.660 519.240 490.920 ;
        RECT 518.520 53.080 518.780 53.340 ;
        RECT 1401.260 53.080 1401.520 53.340 ;
        RECT 1401.260 19.420 1401.520 19.680 ;
        RECT 1407.240 19.420 1407.500 19.680 ;
      LAYER met2 ;
        RECT 520.150 500.000 520.430 504.000 ;
        RECT 520.190 499.790 520.330 500.000 ;
        RECT 520.130 499.470 520.390 499.790 ;
        RECT 518.980 497.090 519.240 497.410 ;
        RECT 519.040 490.950 519.180 497.090 ;
        RECT 518.060 490.630 518.320 490.950 ;
        RECT 518.980 490.630 519.240 490.950 ;
        RECT 518.120 479.640 518.260 490.630 ;
        RECT 518.120 479.500 518.720 479.640 ;
        RECT 518.580 53.370 518.720 479.500 ;
        RECT 518.520 53.050 518.780 53.370 ;
        RECT 1401.260 53.050 1401.520 53.370 ;
        RECT 1401.320 19.710 1401.460 53.050 ;
        RECT 1401.260 19.390 1401.520 19.710 ;
        RECT 1407.240 19.390 1407.500 19.710 ;
        RECT 1407.300 2.400 1407.440 19.390 ;
        RECT 1407.090 -4.800 1407.650 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 478.960 518.350 479.020 ;
        RECT 521.710 478.960 522.030 479.020 ;
        RECT 518.030 478.820 522.030 478.960 ;
        RECT 518.030 478.760 518.350 478.820 ;
        RECT 521.710 478.760 522.030 478.820 ;
        RECT 518.030 52.940 518.350 53.000 ;
        RECT 1423.770 52.940 1424.090 53.000 ;
        RECT 518.030 52.800 1424.090 52.940 ;
        RECT 518.030 52.740 518.350 52.800 ;
        RECT 1423.770 52.740 1424.090 52.800 ;
      LAYER via ;
        RECT 518.060 478.760 518.320 479.020 ;
        RECT 521.740 478.760 522.000 479.020 ;
        RECT 518.060 52.740 518.320 53.000 ;
        RECT 1423.800 52.740 1424.060 53.000 ;
      LAYER met2 ;
        RECT 521.530 500.000 521.810 504.000 ;
        RECT 521.570 498.680 521.710 500.000 ;
        RECT 521.570 498.540 521.940 498.680 ;
        RECT 521.800 479.050 521.940 498.540 ;
        RECT 518.060 478.730 518.320 479.050 ;
        RECT 521.740 478.730 522.000 479.050 ;
        RECT 518.120 53.030 518.260 478.730 ;
        RECT 518.060 52.710 518.320 53.030 ;
        RECT 1423.800 52.710 1424.060 53.030 ;
        RECT 1423.860 2.400 1424.000 52.710 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.630 445.980 522.950 446.040 ;
        RECT 1435.270 445.980 1435.590 446.040 ;
        RECT 522.630 445.840 1435.590 445.980 ;
        RECT 522.630 445.780 522.950 445.840 ;
        RECT 1435.270 445.780 1435.590 445.840 ;
      LAYER via ;
        RECT 522.660 445.780 522.920 446.040 ;
        RECT 1435.300 445.780 1435.560 446.040 ;
      LAYER met2 ;
        RECT 522.910 500.000 523.190 504.000 ;
        RECT 522.950 499.645 523.090 500.000 ;
        RECT 522.880 499.275 523.160 499.645 ;
        RECT 522.650 497.915 522.930 498.285 ;
        RECT 522.720 446.070 522.860 497.915 ;
        RECT 522.660 445.750 522.920 446.070 ;
        RECT 1435.300 445.750 1435.560 446.070 ;
        RECT 1435.360 82.870 1435.500 445.750 ;
        RECT 1435.360 82.730 1440.560 82.870 ;
        RECT 1440.420 2.400 1440.560 82.730 ;
        RECT 1440.210 -4.800 1440.770 2.400 ;
      LAYER via2 ;
        RECT 522.880 499.320 523.160 499.600 ;
        RECT 522.650 497.960 522.930 498.240 ;
      LAYER met3 ;
        RECT 522.855 499.295 523.185 499.625 ;
        RECT 522.870 498.265 523.170 499.295 ;
        RECT 522.625 497.950 523.170 498.265 ;
        RECT 522.625 497.935 522.955 497.950 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.240 500.180 524.560 500.440 ;
        RECT 524.330 499.700 524.470 500.180 ;
        RECT 524.330 499.560 524.700 499.700 ;
        RECT 524.560 498.740 524.700 499.560 ;
        RECT 524.470 498.480 524.790 498.740 ;
        RECT 524.470 487.800 524.790 487.860 ;
        RECT 569.090 487.800 569.410 487.860 ;
        RECT 524.470 487.660 569.410 487.800 ;
        RECT 524.470 487.600 524.790 487.660 ;
        RECT 569.090 487.600 569.410 487.660 ;
        RECT 569.090 483.720 569.410 483.780 ;
        RECT 598.530 483.720 598.850 483.780 ;
        RECT 569.090 483.580 598.850 483.720 ;
        RECT 569.090 483.520 569.410 483.580 ;
        RECT 598.530 483.520 598.850 483.580 ;
        RECT 598.530 452.780 598.850 452.840 ;
        RECT 1455.970 452.780 1456.290 452.840 ;
        RECT 598.530 452.640 1456.290 452.780 ;
        RECT 598.530 452.580 598.850 452.640 ;
        RECT 1455.970 452.580 1456.290 452.640 ;
      LAYER via ;
        RECT 524.270 500.180 524.530 500.440 ;
        RECT 524.500 498.480 524.760 498.740 ;
        RECT 524.500 487.600 524.760 487.860 ;
        RECT 569.120 487.600 569.380 487.860 ;
        RECT 569.120 483.520 569.380 483.780 ;
        RECT 598.560 483.520 598.820 483.780 ;
        RECT 598.560 452.580 598.820 452.840 ;
        RECT 1456.000 452.580 1456.260 452.840 ;
      LAYER met2 ;
        RECT 524.290 500.470 524.570 504.000 ;
        RECT 524.270 500.150 524.570 500.470 ;
        RECT 524.290 500.000 524.570 500.150 ;
        RECT 524.500 498.450 524.760 498.770 ;
        RECT 524.560 487.890 524.700 498.450 ;
        RECT 524.500 487.570 524.760 487.890 ;
        RECT 569.120 487.570 569.380 487.890 ;
        RECT 569.180 483.810 569.320 487.570 ;
        RECT 569.120 483.490 569.380 483.810 ;
        RECT 598.560 483.490 598.820 483.810 ;
        RECT 598.620 452.870 598.760 483.490 ;
        RECT 598.560 452.550 598.820 452.870 ;
        RECT 1456.000 452.550 1456.260 452.870 ;
        RECT 1456.060 17.410 1456.200 452.550 ;
        RECT 1456.060 17.270 1457.120 17.410 ;
        RECT 1456.980 2.400 1457.120 17.270 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.620 499.500 525.940 499.760 ;
        RECT 525.710 498.060 525.850 499.500 ;
        RECT 525.390 497.860 525.850 498.060 ;
        RECT 525.390 497.800 525.710 497.860 ;
        RECT 525.390 479.980 525.710 480.040 ;
        RECT 528.610 479.980 528.930 480.040 ;
        RECT 525.390 479.840 528.930 479.980 ;
        RECT 525.390 479.780 525.710 479.840 ;
        RECT 528.610 479.780 528.930 479.840 ;
        RECT 528.610 445.640 528.930 445.700 ;
        RECT 1469.770 445.640 1470.090 445.700 ;
        RECT 528.610 445.500 1470.090 445.640 ;
        RECT 528.610 445.440 528.930 445.500 ;
        RECT 1469.770 445.440 1470.090 445.500 ;
      LAYER via ;
        RECT 525.650 499.500 525.910 499.760 ;
        RECT 525.420 497.800 525.680 498.060 ;
        RECT 525.420 479.780 525.680 480.040 ;
        RECT 528.640 479.780 528.900 480.040 ;
        RECT 528.640 445.440 528.900 445.700 ;
        RECT 1469.800 445.440 1470.060 445.700 ;
      LAYER met2 ;
        RECT 525.670 500.000 525.950 504.000 ;
        RECT 525.710 499.790 525.850 500.000 ;
        RECT 525.650 499.470 525.910 499.790 ;
        RECT 525.420 497.770 525.680 498.090 ;
        RECT 525.480 480.070 525.620 497.770 ;
        RECT 525.420 479.750 525.680 480.070 ;
        RECT 528.640 479.750 528.900 480.070 ;
        RECT 528.700 445.730 528.840 479.750 ;
        RECT 528.640 445.410 528.900 445.730 ;
        RECT 1469.800 445.410 1470.060 445.730 ;
        RECT 1469.860 82.870 1470.000 445.410 ;
        RECT 1469.860 82.730 1473.680 82.870 ;
        RECT 1473.540 2.400 1473.680 82.730 ;
        RECT 1473.330 -4.800 1473.890 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.000 499.160 527.320 499.420 ;
        RECT 527.090 497.720 527.230 499.160 ;
        RECT 527.090 497.520 527.550 497.720 ;
        RECT 527.230 497.460 527.550 497.520 ;
        RECT 525.390 479.300 525.710 479.360 ;
        RECT 526.770 479.300 527.090 479.360 ;
        RECT 525.390 479.160 527.090 479.300 ;
        RECT 525.390 479.100 525.710 479.160 ;
        RECT 526.770 479.100 527.090 479.160 ;
        RECT 525.390 52.600 525.710 52.660 ;
        RECT 1484.030 52.600 1484.350 52.660 ;
        RECT 525.390 52.460 1484.350 52.600 ;
        RECT 525.390 52.400 525.710 52.460 ;
        RECT 1484.030 52.400 1484.350 52.460 ;
        RECT 1484.030 20.300 1484.350 20.360 ;
        RECT 1490.010 20.300 1490.330 20.360 ;
        RECT 1484.030 20.160 1490.330 20.300 ;
        RECT 1484.030 20.100 1484.350 20.160 ;
        RECT 1490.010 20.100 1490.330 20.160 ;
      LAYER via ;
        RECT 527.030 499.160 527.290 499.420 ;
        RECT 527.260 497.460 527.520 497.720 ;
        RECT 525.420 479.100 525.680 479.360 ;
        RECT 526.800 479.100 527.060 479.360 ;
        RECT 525.420 52.400 525.680 52.660 ;
        RECT 1484.060 52.400 1484.320 52.660 ;
        RECT 1484.060 20.100 1484.320 20.360 ;
        RECT 1490.040 20.100 1490.300 20.360 ;
      LAYER met2 ;
        RECT 527.050 500.000 527.330 504.000 ;
        RECT 527.090 499.450 527.230 500.000 ;
        RECT 527.030 499.130 527.290 499.450 ;
        RECT 527.260 497.660 527.520 497.750 ;
        RECT 526.860 497.520 527.520 497.660 ;
        RECT 526.860 479.390 527.000 497.520 ;
        RECT 527.260 497.430 527.520 497.520 ;
        RECT 525.420 479.070 525.680 479.390 ;
        RECT 526.800 479.070 527.060 479.390 ;
        RECT 525.480 52.690 525.620 479.070 ;
        RECT 525.420 52.370 525.680 52.690 ;
        RECT 1484.060 52.370 1484.320 52.690 ;
        RECT 1484.120 20.390 1484.260 52.370 ;
        RECT 1484.060 20.070 1484.320 20.390 ;
        RECT 1490.040 20.070 1490.300 20.390 ;
        RECT 1490.100 2.400 1490.240 20.070 ;
        RECT 1489.890 -4.800 1490.450 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.850 484.400 526.170 484.460 ;
        RECT 528.150 484.400 528.470 484.460 ;
        RECT 525.850 484.260 528.470 484.400 ;
        RECT 525.850 484.200 526.170 484.260 ;
        RECT 528.150 484.200 528.470 484.260 ;
        RECT 524.930 477.940 525.250 478.000 ;
        RECT 525.850 477.940 526.170 478.000 ;
        RECT 524.930 477.800 526.170 477.940 ;
        RECT 524.930 477.740 525.250 477.800 ;
        RECT 525.850 477.740 526.170 477.800 ;
        RECT 524.930 52.260 525.250 52.320 ;
        RECT 1506.570 52.260 1506.890 52.320 ;
        RECT 524.930 52.120 1506.890 52.260 ;
        RECT 524.930 52.060 525.250 52.120 ;
        RECT 1506.570 52.060 1506.890 52.120 ;
      LAYER via ;
        RECT 525.880 484.200 526.140 484.460 ;
        RECT 528.180 484.200 528.440 484.460 ;
        RECT 524.960 477.740 525.220 478.000 ;
        RECT 525.880 477.740 526.140 478.000 ;
        RECT 524.960 52.060 525.220 52.320 ;
        RECT 1506.600 52.060 1506.860 52.320 ;
      LAYER met2 ;
        RECT 528.430 500.000 528.710 504.000 ;
        RECT 528.470 498.680 528.610 500.000 ;
        RECT 528.240 498.540 528.610 498.680 ;
        RECT 528.240 484.490 528.380 498.540 ;
        RECT 525.880 484.170 526.140 484.490 ;
        RECT 528.180 484.170 528.440 484.490 ;
        RECT 525.940 478.030 526.080 484.170 ;
        RECT 524.960 477.710 525.220 478.030 ;
        RECT 525.880 477.710 526.140 478.030 ;
        RECT 525.020 52.350 525.160 477.710 ;
        RECT 524.960 52.030 525.220 52.350 ;
        RECT 1506.600 52.030 1506.860 52.350 ;
        RECT 1506.660 2.400 1506.800 52.030 ;
        RECT 1506.450 -4.800 1507.010 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.250 748.580 406.570 748.640 ;
        RECT 445.810 748.580 446.130 748.640 ;
        RECT 406.250 748.440 446.130 748.580 ;
        RECT 406.250 748.380 406.570 748.440 ;
        RECT 445.810 748.380 446.130 748.440 ;
        RECT 466.280 499.500 466.600 499.760 ;
        RECT 466.370 499.360 466.510 499.500 ;
        RECT 466.140 499.220 466.510 499.360 ;
        RECT 466.140 498.060 466.280 499.220 ;
        RECT 466.050 497.800 466.370 498.060 ;
        RECT 406.250 480.320 406.570 480.380 ;
        RECT 466.050 480.320 466.370 480.380 ;
        RECT 406.250 480.180 466.370 480.320 ;
        RECT 406.250 480.120 406.570 480.180 ;
        RECT 466.050 480.120 466.370 480.180 ;
        RECT 466.050 61.100 466.370 61.160 ;
        RECT 761.370 61.100 761.690 61.160 ;
        RECT 466.050 60.960 761.690 61.100 ;
        RECT 466.050 60.900 466.370 60.960 ;
        RECT 761.370 60.900 761.690 60.960 ;
      LAYER via ;
        RECT 406.280 748.380 406.540 748.640 ;
        RECT 445.840 748.380 446.100 748.640 ;
        RECT 466.310 499.500 466.570 499.760 ;
        RECT 466.080 497.800 466.340 498.060 ;
        RECT 406.280 480.120 406.540 480.380 ;
        RECT 466.080 480.120 466.340 480.380 ;
        RECT 466.080 60.900 466.340 61.160 ;
        RECT 761.400 60.900 761.660 61.160 ;
      LAYER met2 ;
        RECT 406.280 748.350 406.540 748.670 ;
        RECT 445.840 748.410 446.100 748.670 ;
        RECT 446.550 748.410 446.830 750.000 ;
        RECT 445.840 748.350 446.830 748.410 ;
        RECT 406.340 480.410 406.480 748.350 ;
        RECT 445.900 748.270 446.830 748.350 ;
        RECT 446.550 746.000 446.830 748.270 ;
        RECT 466.330 500.000 466.610 504.000 ;
        RECT 466.370 499.790 466.510 500.000 ;
        RECT 466.310 499.470 466.570 499.790 ;
        RECT 466.080 497.770 466.340 498.090 ;
        RECT 466.140 480.410 466.280 497.770 ;
        RECT 406.280 480.090 406.540 480.410 ;
        RECT 466.080 480.090 466.340 480.410 ;
        RECT 466.140 61.190 466.280 480.090 ;
        RECT 466.080 60.870 466.340 61.190 ;
        RECT 761.400 60.870 761.660 61.190 ;
        RECT 761.460 2.400 761.600 60.870 ;
        RECT 761.250 -4.800 761.810 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 529.760 499.360 530.080 499.420 ;
        RECT 529.760 499.160 530.220 499.360 ;
        RECT 530.080 498.740 530.220 499.160 ;
        RECT 529.990 498.480 530.310 498.740 ;
        RECT 525.850 469.780 526.170 469.840 ;
        RECT 529.530 469.780 529.850 469.840 ;
        RECT 525.850 469.640 529.850 469.780 ;
        RECT 525.850 469.580 526.170 469.640 ;
        RECT 529.530 469.580 529.850 469.640 ;
        RECT 525.850 51.920 526.170 51.980 ;
        RECT 1523.130 51.920 1523.450 51.980 ;
        RECT 525.850 51.780 1523.450 51.920 ;
        RECT 525.850 51.720 526.170 51.780 ;
        RECT 1523.130 51.720 1523.450 51.780 ;
      LAYER via ;
        RECT 529.790 499.160 530.050 499.420 ;
        RECT 530.020 498.480 530.280 498.740 ;
        RECT 525.880 469.580 526.140 469.840 ;
        RECT 529.560 469.580 529.820 469.840 ;
        RECT 525.880 51.720 526.140 51.980 ;
        RECT 1523.160 51.720 1523.420 51.980 ;
      LAYER met2 ;
        RECT 529.810 500.000 530.090 504.000 ;
        RECT 529.850 499.450 529.990 500.000 ;
        RECT 529.790 499.130 530.050 499.450 ;
        RECT 530.020 498.450 530.280 498.770 ;
        RECT 530.080 497.490 530.220 498.450 ;
        RECT 529.620 497.350 530.220 497.490 ;
        RECT 529.620 469.870 529.760 497.350 ;
        RECT 525.880 469.550 526.140 469.870 ;
        RECT 529.560 469.550 529.820 469.870 ;
        RECT 525.940 52.010 526.080 469.550 ;
        RECT 525.880 51.690 526.140 52.010 ;
        RECT 1523.160 51.690 1523.420 52.010 ;
        RECT 1523.220 2.400 1523.360 51.690 ;
        RECT 1523.010 -4.800 1523.570 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.140 499.500 531.460 499.760 ;
        RECT 531.230 499.020 531.370 499.500 ;
        RECT 531.000 498.880 531.370 499.020 ;
        RECT 531.000 498.400 531.140 498.880 ;
        RECT 530.910 498.140 531.230 498.400 ;
        RECT 530.910 487.460 531.230 487.520 ;
        RECT 569.550 487.460 569.870 487.520 ;
        RECT 530.910 487.320 569.870 487.460 ;
        RECT 530.910 487.260 531.230 487.320 ;
        RECT 569.550 487.260 569.870 487.320 ;
        RECT 569.550 452.440 569.870 452.500 ;
        RECT 1538.770 452.440 1539.090 452.500 ;
        RECT 569.550 452.300 1539.090 452.440 ;
        RECT 569.550 452.240 569.870 452.300 ;
        RECT 1538.770 452.240 1539.090 452.300 ;
      LAYER via ;
        RECT 531.170 499.500 531.430 499.760 ;
        RECT 530.940 498.140 531.200 498.400 ;
        RECT 530.940 487.260 531.200 487.520 ;
        RECT 569.580 487.260 569.840 487.520 ;
        RECT 569.580 452.240 569.840 452.500 ;
        RECT 1538.800 452.240 1539.060 452.500 ;
      LAYER met2 ;
        RECT 531.190 500.000 531.470 504.000 ;
        RECT 531.230 499.790 531.370 500.000 ;
        RECT 531.170 499.470 531.430 499.790 ;
        RECT 530.940 498.110 531.200 498.430 ;
        RECT 531.000 487.550 531.140 498.110 ;
        RECT 530.940 487.230 531.200 487.550 ;
        RECT 569.580 487.230 569.840 487.550 ;
        RECT 569.640 452.530 569.780 487.230 ;
        RECT 569.580 452.210 569.840 452.530 ;
        RECT 1538.800 452.210 1539.060 452.530 ;
        RECT 1538.860 17.410 1539.000 452.210 ;
        RECT 1538.860 17.270 1539.920 17.410 ;
        RECT 1539.780 2.400 1539.920 17.270 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.520 499.500 532.840 499.760 ;
        RECT 532.610 497.380 532.750 499.500 ;
        RECT 532.290 497.180 532.750 497.380 ;
        RECT 532.290 497.120 532.610 497.180 ;
        RECT 532.290 483.720 532.610 483.780 ;
        RECT 535.510 483.720 535.830 483.780 ;
        RECT 532.290 483.580 535.830 483.720 ;
        RECT 532.290 483.520 532.610 483.580 ;
        RECT 535.510 483.520 535.830 483.580 ;
        RECT 535.510 452.100 535.830 452.160 ;
        RECT 1552.570 452.100 1552.890 452.160 ;
        RECT 535.510 451.960 1552.890 452.100 ;
        RECT 535.510 451.900 535.830 451.960 ;
        RECT 1552.570 451.900 1552.890 451.960 ;
      LAYER via ;
        RECT 532.550 499.500 532.810 499.760 ;
        RECT 532.320 497.120 532.580 497.380 ;
        RECT 532.320 483.520 532.580 483.780 ;
        RECT 535.540 483.520 535.800 483.780 ;
        RECT 535.540 451.900 535.800 452.160 ;
        RECT 1552.600 451.900 1552.860 452.160 ;
      LAYER met2 ;
        RECT 532.570 500.000 532.850 504.000 ;
        RECT 532.610 499.790 532.750 500.000 ;
        RECT 532.550 499.470 532.810 499.790 ;
        RECT 532.320 497.090 532.580 497.410 ;
        RECT 532.380 483.810 532.520 497.090 ;
        RECT 532.320 483.490 532.580 483.810 ;
        RECT 535.540 483.490 535.800 483.810 ;
        RECT 535.600 452.190 535.740 483.490 ;
        RECT 535.540 451.870 535.800 452.190 ;
        RECT 1552.600 451.870 1552.860 452.190 ;
        RECT 1552.660 82.870 1552.800 451.870 ;
        RECT 1552.660 82.730 1556.480 82.870 ;
        RECT 1556.340 2.400 1556.480 82.730 ;
        RECT 1556.130 -4.800 1556.690 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.130 480.660 534.450 480.720 ;
        RECT 534.130 480.520 535.740 480.660 ;
        RECT 534.130 480.460 534.450 480.520 ;
        RECT 535.050 479.640 535.370 479.700 ;
        RECT 535.600 479.640 535.740 480.520 ;
        RECT 535.050 479.500 535.740 479.640 ;
        RECT 535.050 479.440 535.370 479.500 ;
        RECT 535.050 411.300 535.370 411.360 ;
        RECT 1566.370 411.300 1566.690 411.360 ;
        RECT 535.050 411.160 1566.690 411.300 ;
        RECT 535.050 411.100 535.370 411.160 ;
        RECT 1566.370 411.100 1566.690 411.160 ;
        RECT 1566.370 16.900 1566.690 16.960 ;
        RECT 1572.810 16.900 1573.130 16.960 ;
        RECT 1566.370 16.760 1573.130 16.900 ;
        RECT 1566.370 16.700 1566.690 16.760 ;
        RECT 1572.810 16.700 1573.130 16.760 ;
      LAYER via ;
        RECT 534.160 480.460 534.420 480.720 ;
        RECT 535.080 479.440 535.340 479.700 ;
        RECT 535.080 411.100 535.340 411.360 ;
        RECT 1566.400 411.100 1566.660 411.360 ;
        RECT 1566.400 16.700 1566.660 16.960 ;
        RECT 1572.840 16.700 1573.100 16.960 ;
      LAYER met2 ;
        RECT 533.950 500.000 534.230 504.000 ;
        RECT 533.990 498.680 534.130 500.000 ;
        RECT 533.990 498.540 534.360 498.680 ;
        RECT 534.220 480.750 534.360 498.540 ;
        RECT 534.160 480.430 534.420 480.750 ;
        RECT 535.080 479.410 535.340 479.730 ;
        RECT 535.140 411.390 535.280 479.410 ;
        RECT 535.080 411.070 535.340 411.390 ;
        RECT 1566.400 411.070 1566.660 411.390 ;
        RECT 1566.460 16.990 1566.600 411.070 ;
        RECT 1566.400 16.670 1566.660 16.990 ;
        RECT 1572.840 16.670 1573.100 16.990 ;
        RECT 1572.900 2.400 1573.040 16.670 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.280 499.500 535.600 499.760 ;
        RECT 535.370 498.740 535.510 499.500 ;
        RECT 535.050 498.540 535.510 498.740 ;
        RECT 535.050 498.480 535.370 498.540 ;
        RECT 531.830 480.320 532.150 480.380 ;
        RECT 535.050 480.320 535.370 480.380 ;
        RECT 531.830 480.180 535.370 480.320 ;
        RECT 531.830 480.120 532.150 480.180 ;
        RECT 535.050 480.120 535.370 480.180 ;
        RECT 531.830 60.760 532.150 60.820 ;
        RECT 1589.370 60.760 1589.690 60.820 ;
        RECT 531.830 60.620 1589.690 60.760 ;
        RECT 531.830 60.560 532.150 60.620 ;
        RECT 1589.370 60.560 1589.690 60.620 ;
      LAYER via ;
        RECT 535.310 499.500 535.570 499.760 ;
        RECT 535.080 498.480 535.340 498.740 ;
        RECT 531.860 480.120 532.120 480.380 ;
        RECT 535.080 480.120 535.340 480.380 ;
        RECT 531.860 60.560 532.120 60.820 ;
        RECT 1589.400 60.560 1589.660 60.820 ;
      LAYER met2 ;
        RECT 535.330 500.000 535.610 504.000 ;
        RECT 535.370 499.790 535.510 500.000 ;
        RECT 535.310 499.470 535.570 499.790 ;
        RECT 535.080 498.450 535.340 498.770 ;
        RECT 535.140 480.410 535.280 498.450 ;
        RECT 531.860 480.090 532.120 480.410 ;
        RECT 535.080 480.090 535.340 480.410 ;
        RECT 531.920 60.850 532.060 480.090 ;
        RECT 531.860 60.530 532.120 60.850 ;
        RECT 1589.400 60.530 1589.660 60.850 ;
        RECT 1589.460 2.400 1589.600 60.530 ;
        RECT 1589.250 -4.800 1589.810 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 536.660 500.180 536.980 500.440 ;
        RECT 536.750 499.700 536.890 500.180 ;
        RECT 536.750 499.560 537.580 499.700 ;
        RECT 537.440 498.740 537.580 499.560 ;
        RECT 537.350 498.480 537.670 498.740 ;
      LAYER via ;
        RECT 536.690 500.180 536.950 500.440 ;
        RECT 537.380 498.480 537.640 498.740 ;
      LAYER met2 ;
        RECT 536.710 500.470 536.990 504.000 ;
        RECT 536.690 500.150 536.990 500.470 ;
        RECT 536.710 500.000 536.990 500.150 ;
        RECT 537.380 498.450 537.640 498.770 ;
        RECT 537.440 498.285 537.580 498.450 ;
        RECT 537.370 497.915 537.650 498.285 ;
        RECT 1605.950 57.955 1606.230 58.325 ;
        RECT 1606.020 2.400 1606.160 57.955 ;
        RECT 1605.810 -4.800 1606.370 2.400 ;
      LAYER via2 ;
        RECT 537.370 497.960 537.650 498.240 ;
        RECT 1605.950 58.000 1606.230 58.280 ;
      LAYER met3 ;
        RECT 537.345 498.260 537.675 498.265 ;
        RECT 537.345 498.250 537.930 498.260 ;
        RECT 537.345 497.950 538.130 498.250 ;
        RECT 537.345 497.940 537.930 497.950 ;
        RECT 537.345 497.935 537.675 497.940 ;
        RECT 537.550 58.290 537.930 58.300 ;
        RECT 1605.925 58.290 1606.255 58.305 ;
        RECT 537.550 57.990 1606.255 58.290 ;
        RECT 537.550 57.980 537.930 57.990 ;
        RECT 1605.925 57.975 1606.255 57.990 ;
      LAYER via3 ;
        RECT 537.580 497.940 537.900 498.260 ;
        RECT 537.580 57.980 537.900 58.300 ;
      LAYER met4 ;
        RECT 537.575 497.935 537.905 498.265 ;
        RECT 537.590 58.305 537.890 497.935 ;
        RECT 537.575 57.975 537.905 58.305 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.040 499.500 538.360 499.760 ;
        RECT 538.130 499.080 538.270 499.500 ;
        RECT 538.130 498.880 538.590 499.080 ;
        RECT 538.270 498.820 538.590 498.880 ;
        RECT 538.730 477.940 539.050 478.000 ;
        RECT 543.790 477.940 544.110 478.000 ;
        RECT 538.730 477.800 544.110 477.940 ;
        RECT 538.730 477.740 539.050 477.800 ;
        RECT 543.790 477.740 544.110 477.800 ;
        RECT 543.790 425.580 544.110 425.640 ;
        RECT 1621.570 425.580 1621.890 425.640 ;
        RECT 543.790 425.440 1621.890 425.580 ;
        RECT 543.790 425.380 544.110 425.440 ;
        RECT 1621.570 425.380 1621.890 425.440 ;
      LAYER via ;
        RECT 538.070 499.500 538.330 499.760 ;
        RECT 538.300 498.820 538.560 499.080 ;
        RECT 538.760 477.740 539.020 478.000 ;
        RECT 543.820 477.740 544.080 478.000 ;
        RECT 543.820 425.380 544.080 425.640 ;
        RECT 1621.600 425.380 1621.860 425.640 ;
      LAYER met2 ;
        RECT 538.090 500.000 538.370 504.000 ;
        RECT 538.130 499.790 538.270 500.000 ;
        RECT 538.070 499.470 538.330 499.790 ;
        RECT 538.300 498.790 538.560 499.110 ;
        RECT 538.360 498.340 538.500 498.790 ;
        RECT 538.360 498.200 538.960 498.340 ;
        RECT 538.820 478.030 538.960 498.200 ;
        RECT 538.760 477.710 539.020 478.030 ;
        RECT 543.820 477.710 544.080 478.030 ;
        RECT 543.880 425.670 544.020 477.710 ;
        RECT 543.820 425.350 544.080 425.670 ;
        RECT 1621.600 425.350 1621.860 425.670 ;
        RECT 1621.660 17.410 1621.800 425.350 ;
        RECT 1621.660 17.270 1622.720 17.410 ;
        RECT 1622.580 2.400 1622.720 17.270 ;
        RECT 1622.370 -4.800 1622.930 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 60.080 538.590 60.140 ;
        RECT 1639.050 60.080 1639.370 60.140 ;
        RECT 538.270 59.940 1639.370 60.080 ;
        RECT 538.270 59.880 538.590 59.940 ;
        RECT 1639.050 59.880 1639.370 59.940 ;
      LAYER via ;
        RECT 538.300 59.880 538.560 60.140 ;
        RECT 1639.080 59.880 1639.340 60.140 ;
      LAYER met2 ;
        RECT 539.470 500.000 539.750 504.000 ;
        RECT 539.510 499.815 539.650 500.000 ;
        RECT 539.440 499.445 539.720 499.815 ;
        RECT 538.290 497.235 538.570 497.605 ;
        RECT 538.360 60.170 538.500 497.235 ;
        RECT 538.300 59.850 538.560 60.170 ;
        RECT 1639.080 59.850 1639.340 60.170 ;
        RECT 1639.140 2.400 1639.280 59.850 ;
        RECT 1638.930 -4.800 1639.490 2.400 ;
      LAYER via2 ;
        RECT 539.440 499.490 539.720 499.770 ;
        RECT 538.290 497.280 538.570 497.560 ;
      LAYER met3 ;
        RECT 539.415 499.465 539.745 499.795 ;
        RECT 538.265 497.570 538.595 497.585 ;
        RECT 539.430 497.570 539.730 499.465 ;
        RECT 538.265 497.270 539.730 497.570 ;
        RECT 538.265 497.255 538.595 497.270 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 470.120 539.510 470.180 ;
        RECT 541.030 470.120 541.350 470.180 ;
        RECT 539.190 469.980 541.350 470.120 ;
        RECT 539.190 469.920 539.510 469.980 ;
        RECT 541.030 469.920 541.350 469.980 ;
        RECT 539.190 59.740 539.510 59.800 ;
        RECT 1649.630 59.740 1649.950 59.800 ;
        RECT 539.190 59.600 1649.950 59.740 ;
        RECT 539.190 59.540 539.510 59.600 ;
        RECT 1649.630 59.540 1649.950 59.600 ;
        RECT 1649.630 20.300 1649.950 20.360 ;
        RECT 1655.610 20.300 1655.930 20.360 ;
        RECT 1649.630 20.160 1655.930 20.300 ;
        RECT 1649.630 20.100 1649.950 20.160 ;
        RECT 1655.610 20.100 1655.930 20.160 ;
      LAYER via ;
        RECT 539.220 469.920 539.480 470.180 ;
        RECT 541.060 469.920 541.320 470.180 ;
        RECT 539.220 59.540 539.480 59.800 ;
        RECT 1649.660 59.540 1649.920 59.800 ;
        RECT 1649.660 20.100 1649.920 20.360 ;
        RECT 1655.640 20.100 1655.900 20.360 ;
      LAYER met2 ;
        RECT 540.850 500.000 541.130 504.000 ;
        RECT 540.890 498.680 541.030 500.000 ;
        RECT 540.890 498.540 541.260 498.680 ;
        RECT 541.120 470.210 541.260 498.540 ;
        RECT 539.220 469.890 539.480 470.210 ;
        RECT 541.060 469.890 541.320 470.210 ;
        RECT 539.280 59.830 539.420 469.890 ;
        RECT 539.220 59.510 539.480 59.830 ;
        RECT 1649.660 59.510 1649.920 59.830 ;
        RECT 1649.720 20.390 1649.860 59.510 ;
        RECT 1649.660 20.070 1649.920 20.390 ;
        RECT 1655.640 20.070 1655.900 20.390 ;
        RECT 1655.700 2.400 1655.840 20.070 ;
        RECT 1655.490 -4.800 1656.050 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 59.400 539.050 59.460 ;
        RECT 1672.170 59.400 1672.490 59.460 ;
        RECT 538.730 59.260 1672.490 59.400 ;
        RECT 538.730 59.200 539.050 59.260 ;
        RECT 1672.170 59.200 1672.490 59.260 ;
      LAYER via ;
        RECT 538.760 59.200 539.020 59.460 ;
        RECT 1672.200 59.200 1672.460 59.460 ;
      LAYER met2 ;
        RECT 542.230 500.000 542.510 504.000 ;
        RECT 542.270 499.020 542.410 500.000 ;
        RECT 542.040 498.965 542.410 499.020 ;
        RECT 541.970 498.880 542.410 498.965 ;
        RECT 541.970 498.595 542.250 498.880 ;
        RECT 538.750 476.835 539.030 477.205 ;
        RECT 538.820 59.490 538.960 476.835 ;
        RECT 538.760 59.170 539.020 59.490 ;
        RECT 1672.200 59.170 1672.460 59.490 ;
        RECT 1672.260 2.400 1672.400 59.170 ;
        RECT 1672.050 -4.800 1672.610 2.400 ;
      LAYER via2 ;
        RECT 541.970 498.640 542.250 498.920 ;
        RECT 538.750 476.880 539.030 477.160 ;
      LAYER met3 ;
        RECT 540.310 498.930 540.690 498.940 ;
        RECT 541.945 498.930 542.275 498.945 ;
        RECT 540.310 498.630 542.275 498.930 ;
        RECT 540.310 498.620 540.690 498.630 ;
        RECT 541.945 498.615 542.275 498.630 ;
        RECT 538.725 477.170 539.055 477.185 ;
        RECT 540.310 477.170 540.690 477.180 ;
        RECT 538.725 476.870 540.690 477.170 ;
        RECT 538.725 476.855 539.055 476.870 ;
        RECT 540.310 476.860 540.690 476.870 ;
      LAYER via3 ;
        RECT 540.340 498.620 540.660 498.940 ;
        RECT 540.340 476.860 540.660 477.180 ;
      LAYER met4 ;
        RECT 540.335 498.615 540.665 498.945 ;
        RECT 540.350 477.185 540.650 498.615 ;
        RECT 540.335 476.855 540.665 477.185 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 405.790 749.600 406.110 749.660 ;
        RECT 405.790 749.460 446.960 749.600 ;
        RECT 405.790 749.400 406.110 749.460 ;
        RECT 446.820 748.920 446.960 749.460 ;
        RECT 451.330 748.920 451.650 748.980 ;
        RECT 446.820 748.780 451.650 748.920 ;
        RECT 451.330 748.720 451.650 748.780 ;
        RECT 466.510 497.320 466.830 497.380 ;
        RECT 467.890 497.320 468.210 497.380 ;
        RECT 466.510 497.180 468.210 497.320 ;
        RECT 466.510 497.120 466.830 497.180 ;
        RECT 467.890 497.120 468.210 497.180 ;
        RECT 405.790 479.300 406.110 479.360 ;
        RECT 466.510 479.300 466.830 479.360 ;
        RECT 405.790 479.160 466.830 479.300 ;
        RECT 405.790 479.100 406.110 479.160 ;
        RECT 466.510 479.100 466.830 479.160 ;
        RECT 466.510 67.560 466.830 67.620 ;
        RECT 777.930 67.560 778.250 67.620 ;
        RECT 466.510 67.420 778.250 67.560 ;
        RECT 466.510 67.360 466.830 67.420 ;
        RECT 777.930 67.360 778.250 67.420 ;
      LAYER via ;
        RECT 405.820 749.400 406.080 749.660 ;
        RECT 451.360 748.720 451.620 748.980 ;
        RECT 466.540 497.120 466.800 497.380 ;
        RECT 467.920 497.120 468.180 497.380 ;
        RECT 405.820 479.100 406.080 479.360 ;
        RECT 466.540 479.100 466.800 479.360 ;
        RECT 466.540 67.360 466.800 67.620 ;
        RECT 777.960 67.360 778.220 67.620 ;
      LAYER met2 ;
        RECT 405.820 749.370 406.080 749.690 ;
        RECT 405.880 479.390 406.020 749.370 ;
        RECT 452.070 749.090 452.350 750.000 ;
        RECT 451.420 749.010 452.350 749.090 ;
        RECT 451.360 748.950 452.350 749.010 ;
        RECT 451.360 748.690 451.620 748.950 ;
        RECT 452.070 746.000 452.350 748.950 ;
        RECT 467.710 500.000 467.990 504.000 ;
        RECT 467.750 498.680 467.890 500.000 ;
        RECT 467.750 498.540 468.120 498.680 ;
        RECT 467.980 497.410 468.120 498.540 ;
        RECT 466.540 497.090 466.800 497.410 ;
        RECT 467.920 497.090 468.180 497.410 ;
        RECT 466.600 479.390 466.740 497.090 ;
        RECT 405.820 479.070 406.080 479.390 ;
        RECT 466.540 479.070 466.800 479.390 ;
        RECT 466.600 67.650 466.740 479.070 ;
        RECT 466.540 67.330 466.800 67.650 ;
        RECT 777.960 67.330 778.220 67.650 ;
        RECT 778.020 2.400 778.160 67.330 ;
        RECT 777.810 -4.800 778.370 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.610 500.000 543.890 504.000 ;
        RECT 543.650 498.340 543.790 500.000 ;
        RECT 543.420 498.285 543.790 498.340 ;
        RECT 543.350 498.200 543.790 498.285 ;
        RECT 543.350 497.915 543.630 498.200 ;
        RECT 1683.690 196.675 1683.970 197.045 ;
        RECT 1683.760 82.870 1683.900 196.675 ;
        RECT 1683.760 82.730 1688.960 82.870 ;
        RECT 1688.820 2.400 1688.960 82.730 ;
        RECT 1688.610 -4.800 1689.170 2.400 ;
      LAYER via2 ;
        RECT 543.350 497.960 543.630 498.240 ;
        RECT 1683.690 196.720 1683.970 197.000 ;
      LAYER met3 ;
        RECT 542.150 498.250 542.530 498.260 ;
        RECT 543.325 498.250 543.655 498.265 ;
        RECT 542.150 497.950 543.655 498.250 ;
        RECT 542.150 497.940 542.530 497.950 ;
        RECT 543.325 497.935 543.655 497.950 ;
        RECT 542.150 197.010 542.530 197.020 ;
        RECT 1683.665 197.010 1683.995 197.025 ;
        RECT 542.150 196.710 1683.995 197.010 ;
        RECT 542.150 196.700 542.530 196.710 ;
        RECT 1683.665 196.695 1683.995 196.710 ;
      LAYER via3 ;
        RECT 542.180 497.940 542.500 498.260 ;
        RECT 542.180 196.700 542.500 197.020 ;
      LAYER met4 ;
        RECT 542.175 497.935 542.505 498.265 ;
        RECT 542.190 197.025 542.490 497.935 ;
        RECT 542.175 196.695 542.505 197.025 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.940 499.020 545.260 499.080 ;
        RECT 544.800 498.820 545.260 499.020 ;
        RECT 544.800 498.060 544.940 498.820 ;
        RECT 544.710 497.800 545.030 498.060 ;
        RECT 544.250 472.160 544.570 472.220 ;
        RECT 547.930 472.160 548.250 472.220 ;
        RECT 544.250 472.020 548.250 472.160 ;
        RECT 544.250 471.960 544.570 472.020 ;
        RECT 547.930 471.960 548.250 472.020 ;
        RECT 547.930 198.460 548.250 198.520 ;
        RECT 1704.370 198.460 1704.690 198.520 ;
        RECT 547.930 198.320 1704.690 198.460 ;
        RECT 547.930 198.260 548.250 198.320 ;
        RECT 1704.370 198.260 1704.690 198.320 ;
      LAYER via ;
        RECT 544.970 498.820 545.230 499.080 ;
        RECT 544.740 497.800 545.000 498.060 ;
        RECT 544.280 471.960 544.540 472.220 ;
        RECT 547.960 471.960 548.220 472.220 ;
        RECT 547.960 198.260 548.220 198.520 ;
        RECT 1704.400 198.260 1704.660 198.520 ;
      LAYER met2 ;
        RECT 544.990 500.000 545.270 504.000 ;
        RECT 545.030 499.110 545.170 500.000 ;
        RECT 544.970 498.790 545.230 499.110 ;
        RECT 544.740 497.770 545.000 498.090 ;
        RECT 544.800 496.870 544.940 497.770 ;
        RECT 544.340 496.730 544.940 496.870 ;
        RECT 544.340 472.250 544.480 496.730 ;
        RECT 544.280 471.930 544.540 472.250 ;
        RECT 547.960 471.930 548.220 472.250 ;
        RECT 548.020 198.550 548.160 471.930 ;
        RECT 547.960 198.230 548.220 198.550 ;
        RECT 1704.400 198.230 1704.660 198.550 ;
        RECT 1704.460 17.410 1704.600 198.230 ;
        RECT 1704.460 17.270 1705.520 17.410 ;
        RECT 1705.380 2.400 1705.520 17.270 ;
        RECT 1705.170 -4.800 1705.730 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.630 66.540 545.950 66.600 ;
        RECT 1721.850 66.540 1722.170 66.600 ;
        RECT 545.630 66.400 1722.170 66.540 ;
        RECT 545.630 66.340 545.950 66.400 ;
        RECT 1721.850 66.340 1722.170 66.400 ;
      LAYER via ;
        RECT 545.660 66.340 545.920 66.600 ;
        RECT 1721.880 66.340 1722.140 66.600 ;
      LAYER met2 ;
        RECT 546.370 500.000 546.650 504.000 ;
        RECT 546.410 498.850 546.550 500.000 ;
        RECT 546.410 498.710 546.780 498.850 ;
        RECT 546.640 481.170 546.780 498.710 ;
        RECT 545.720 481.030 546.780 481.170 ;
        RECT 545.720 66.630 545.860 481.030 ;
        RECT 545.660 66.310 545.920 66.630 ;
        RECT 1721.880 66.310 1722.140 66.630 ;
        RECT 1721.940 2.400 1722.080 66.310 ;
        RECT 1721.730 -4.800 1722.290 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.550 66.200 546.870 66.260 ;
        RECT 1732.430 66.200 1732.750 66.260 ;
        RECT 546.550 66.060 1732.750 66.200 ;
        RECT 546.550 66.000 546.870 66.060 ;
        RECT 1732.430 66.000 1732.750 66.060 ;
        RECT 1732.430 20.300 1732.750 20.360 ;
        RECT 1738.410 20.300 1738.730 20.360 ;
        RECT 1732.430 20.160 1738.730 20.300 ;
        RECT 1732.430 20.100 1732.750 20.160 ;
        RECT 1738.410 20.100 1738.730 20.160 ;
      LAYER via ;
        RECT 546.580 66.000 546.840 66.260 ;
        RECT 1732.460 66.000 1732.720 66.260 ;
        RECT 1732.460 20.100 1732.720 20.360 ;
        RECT 1738.440 20.100 1738.700 20.360 ;
      LAYER met2 ;
        RECT 547.750 500.000 548.030 504.000 ;
        RECT 547.790 499.020 547.930 500.000 ;
        RECT 547.560 498.880 547.930 499.020 ;
        RECT 547.560 481.170 547.700 498.880 ;
        RECT 547.100 481.030 547.700 481.170 ;
        RECT 547.100 479.810 547.240 481.030 ;
        RECT 546.640 479.670 547.240 479.810 ;
        RECT 546.640 66.290 546.780 479.670 ;
        RECT 546.580 65.970 546.840 66.290 ;
        RECT 1732.460 65.970 1732.720 66.290 ;
        RECT 1732.520 20.390 1732.660 65.970 ;
        RECT 1732.460 20.070 1732.720 20.390 ;
        RECT 1738.440 20.070 1738.700 20.390 ;
        RECT 1738.500 2.400 1738.640 20.070 ;
        RECT 1738.290 -4.800 1738.850 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.080 499.500 549.400 499.760 ;
        RECT 549.170 498.400 549.310 499.500 ;
        RECT 549.170 498.200 549.630 498.400 ;
        RECT 549.310 498.140 549.630 498.200 ;
        RECT 546.090 480.320 546.410 480.380 ;
        RECT 549.310 480.320 549.630 480.380 ;
        RECT 546.090 480.180 549.630 480.320 ;
        RECT 546.090 480.120 546.410 480.180 ;
        RECT 549.310 480.120 549.630 480.180 ;
        RECT 546.090 65.860 546.410 65.920 ;
        RECT 1754.970 65.860 1755.290 65.920 ;
        RECT 546.090 65.720 1755.290 65.860 ;
        RECT 546.090 65.660 546.410 65.720 ;
        RECT 1754.970 65.660 1755.290 65.720 ;
      LAYER via ;
        RECT 549.110 499.500 549.370 499.760 ;
        RECT 549.340 498.140 549.600 498.400 ;
        RECT 546.120 480.120 546.380 480.380 ;
        RECT 549.340 480.120 549.600 480.380 ;
        RECT 546.120 65.660 546.380 65.920 ;
        RECT 1755.000 65.660 1755.260 65.920 ;
      LAYER met2 ;
        RECT 549.130 500.000 549.410 504.000 ;
        RECT 549.170 499.790 549.310 500.000 ;
        RECT 549.110 499.470 549.370 499.790 ;
        RECT 549.340 498.110 549.600 498.430 ;
        RECT 549.400 480.410 549.540 498.110 ;
        RECT 546.120 480.090 546.380 480.410 ;
        RECT 549.340 480.090 549.600 480.410 ;
        RECT 546.180 65.950 546.320 480.090 ;
        RECT 546.120 65.630 546.380 65.950 ;
        RECT 1755.000 65.630 1755.260 65.950 ;
        RECT 1755.060 2.400 1755.200 65.630 ;
        RECT 1754.850 -4.800 1755.410 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.460 499.500 550.780 499.760 ;
        RECT 550.550 499.020 550.690 499.500 ;
        RECT 550.320 498.880 550.690 499.020 ;
        RECT 550.320 498.740 550.460 498.880 ;
        RECT 550.230 498.480 550.550 498.740 ;
      LAYER via ;
        RECT 550.490 499.500 550.750 499.760 ;
        RECT 550.260 498.480 550.520 498.740 ;
      LAYER met2 ;
        RECT 550.510 500.000 550.790 504.000 ;
        RECT 550.550 499.790 550.690 500.000 ;
        RECT 550.490 499.470 550.750 499.790 ;
        RECT 550.260 498.450 550.520 498.770 ;
        RECT 550.320 481.285 550.460 498.450 ;
        RECT 550.250 480.915 550.530 481.285 ;
        RECT 1771.550 64.755 1771.830 65.125 ;
        RECT 1771.620 2.400 1771.760 64.755 ;
        RECT 1771.410 -4.800 1771.970 2.400 ;
      LAYER via2 ;
        RECT 550.250 480.960 550.530 481.240 ;
        RECT 1771.550 64.800 1771.830 65.080 ;
      LAYER met3 ;
        RECT 547.670 481.250 548.050 481.260 ;
        RECT 550.225 481.250 550.555 481.265 ;
        RECT 547.670 480.950 550.555 481.250 ;
        RECT 547.670 480.940 548.050 480.950 ;
        RECT 550.225 480.935 550.555 480.950 ;
        RECT 547.670 65.090 548.050 65.100 ;
        RECT 1771.525 65.090 1771.855 65.105 ;
        RECT 547.670 64.790 1771.855 65.090 ;
        RECT 547.670 64.780 548.050 64.790 ;
        RECT 1771.525 64.775 1771.855 64.790 ;
      LAYER via3 ;
        RECT 547.700 480.940 548.020 481.260 ;
        RECT 547.700 64.780 548.020 65.100 ;
      LAYER met4 ;
        RECT 547.695 480.935 548.025 481.265 ;
        RECT 547.710 65.105 548.010 480.935 ;
        RECT 547.695 64.775 548.025 65.105 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 551.840 499.360 552.160 499.420 ;
        RECT 551.840 499.160 552.300 499.360 ;
        RECT 552.160 498.740 552.300 499.160 ;
        RECT 552.070 498.480 552.390 498.740 ;
        RECT 552.070 486.440 552.390 486.500 ;
        RECT 552.070 486.300 579.670 486.440 ;
        RECT 552.070 486.240 552.390 486.300 ;
        RECT 579.530 485.080 579.670 486.300 ;
        RECT 605.430 485.080 605.750 485.140 ;
        RECT 579.530 484.940 605.750 485.080 ;
        RECT 605.430 484.880 605.750 484.940 ;
        RECT 605.430 460.260 605.750 460.320 ;
        RECT 1787.170 460.260 1787.490 460.320 ;
        RECT 605.430 460.120 1787.490 460.260 ;
        RECT 605.430 460.060 605.750 460.120 ;
        RECT 1787.170 460.060 1787.490 460.120 ;
      LAYER via ;
        RECT 551.870 499.160 552.130 499.420 ;
        RECT 552.100 498.480 552.360 498.740 ;
        RECT 552.100 486.240 552.360 486.500 ;
        RECT 605.460 484.880 605.720 485.140 ;
        RECT 605.460 460.060 605.720 460.320 ;
        RECT 1787.200 460.060 1787.460 460.320 ;
      LAYER met2 ;
        RECT 551.890 500.000 552.170 504.000 ;
        RECT 551.930 499.450 552.070 500.000 ;
        RECT 551.870 499.130 552.130 499.450 ;
        RECT 552.100 498.450 552.360 498.770 ;
        RECT 552.160 486.530 552.300 498.450 ;
        RECT 552.100 486.210 552.360 486.530 ;
        RECT 605.460 484.850 605.720 485.170 ;
        RECT 605.520 460.350 605.660 484.850 ;
        RECT 605.460 460.030 605.720 460.350 ;
        RECT 1787.200 460.030 1787.460 460.350 ;
        RECT 1787.260 17.410 1787.400 460.030 ;
        RECT 1787.260 17.270 1788.320 17.410 ;
        RECT 1788.180 2.400 1788.320 17.270 ;
        RECT 1787.970 -4.800 1788.530 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.990 485.760 553.310 485.820 ;
        RECT 555.750 485.760 556.070 485.820 ;
        RECT 552.990 485.620 556.070 485.760 ;
        RECT 552.990 485.560 553.310 485.620 ;
        RECT 555.750 485.560 556.070 485.620 ;
        RECT 555.750 440.540 556.070 440.600 ;
        RECT 1800.970 440.540 1801.290 440.600 ;
        RECT 555.750 440.400 1801.290 440.540 ;
        RECT 555.750 440.340 556.070 440.400 ;
        RECT 1800.970 440.340 1801.290 440.400 ;
      LAYER via ;
        RECT 553.020 485.560 553.280 485.820 ;
        RECT 555.780 485.560 556.040 485.820 ;
        RECT 555.780 440.340 556.040 440.600 ;
        RECT 1801.000 440.340 1801.260 440.600 ;
      LAYER met2 ;
        RECT 553.270 500.000 553.550 504.000 ;
        RECT 553.310 498.965 553.450 500.000 ;
        RECT 553.240 498.595 553.520 498.965 ;
        RECT 553.010 497.915 553.290 498.285 ;
        RECT 553.080 485.850 553.220 497.915 ;
        RECT 553.020 485.530 553.280 485.850 ;
        RECT 555.780 485.530 556.040 485.850 ;
        RECT 555.840 440.630 555.980 485.530 ;
        RECT 555.780 440.310 556.040 440.630 ;
        RECT 1801.000 440.310 1801.260 440.630 ;
        RECT 1801.060 82.870 1801.200 440.310 ;
        RECT 1801.060 82.730 1804.880 82.870 ;
        RECT 1804.740 2.400 1804.880 82.730 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
      LAYER via2 ;
        RECT 553.240 498.640 553.520 498.920 ;
        RECT 553.010 497.960 553.290 498.240 ;
      LAYER met3 ;
        RECT 553.215 498.615 553.545 498.945 ;
        RECT 553.230 498.265 553.530 498.615 ;
        RECT 552.985 497.950 553.530 498.265 ;
        RECT 552.985 497.935 553.315 497.950 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.830 490.520 555.150 490.580 ;
        RECT 571.390 490.520 571.710 490.580 ;
        RECT 554.830 490.380 571.710 490.520 ;
        RECT 554.830 490.320 555.150 490.380 ;
        RECT 571.390 490.320 571.710 490.380 ;
        RECT 571.390 459.920 571.710 459.980 ;
        RECT 1814.770 459.920 1815.090 459.980 ;
        RECT 571.390 459.780 1815.090 459.920 ;
        RECT 571.390 459.720 571.710 459.780 ;
        RECT 1814.770 459.720 1815.090 459.780 ;
        RECT 1814.770 16.900 1815.090 16.960 ;
        RECT 1821.210 16.900 1821.530 16.960 ;
        RECT 1814.770 16.760 1821.530 16.900 ;
        RECT 1814.770 16.700 1815.090 16.760 ;
        RECT 1821.210 16.700 1821.530 16.760 ;
      LAYER via ;
        RECT 554.860 490.320 555.120 490.580 ;
        RECT 571.420 490.320 571.680 490.580 ;
        RECT 571.420 459.720 571.680 459.980 ;
        RECT 1814.800 459.720 1815.060 459.980 ;
        RECT 1814.800 16.700 1815.060 16.960 ;
        RECT 1821.240 16.700 1821.500 16.960 ;
      LAYER met2 ;
        RECT 554.650 500.000 554.930 504.000 ;
        RECT 554.690 498.680 554.830 500.000 ;
        RECT 554.690 498.540 555.060 498.680 ;
        RECT 554.920 490.610 555.060 498.540 ;
        RECT 554.860 490.290 555.120 490.610 ;
        RECT 571.420 490.290 571.680 490.610 ;
        RECT 571.480 460.010 571.620 490.290 ;
        RECT 571.420 459.690 571.680 460.010 ;
        RECT 1814.800 459.690 1815.060 460.010 ;
        RECT 1814.860 16.990 1815.000 459.690 ;
        RECT 1814.800 16.670 1815.060 16.990 ;
        RECT 1821.240 16.670 1821.500 16.990 ;
        RECT 1821.300 2.400 1821.440 16.670 ;
        RECT 1821.090 -4.800 1821.650 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 65.520 552.390 65.580 ;
        RECT 1837.770 65.520 1838.090 65.580 ;
        RECT 552.070 65.380 1838.090 65.520 ;
        RECT 552.070 65.320 552.390 65.380 ;
        RECT 1837.770 65.320 1838.090 65.380 ;
      LAYER via ;
        RECT 552.100 65.320 552.360 65.580 ;
        RECT 1837.800 65.320 1838.060 65.580 ;
      LAYER met2 ;
        RECT 556.030 500.000 556.310 504.000 ;
        RECT 556.070 499.645 556.210 500.000 ;
        RECT 556.000 499.275 556.280 499.645 ;
        RECT 552.090 482.275 552.370 482.645 ;
        RECT 552.160 65.610 552.300 482.275 ;
        RECT 552.100 65.290 552.360 65.610 ;
        RECT 1837.800 65.290 1838.060 65.610 ;
        RECT 1837.860 2.400 1838.000 65.290 ;
        RECT 1837.650 -4.800 1838.210 2.400 ;
      LAYER via2 ;
        RECT 556.000 499.320 556.280 499.600 ;
        RECT 552.090 482.320 552.370 482.600 ;
      LAYER met3 ;
        RECT 555.030 499.610 555.410 499.620 ;
        RECT 555.975 499.610 556.305 499.625 ;
        RECT 555.030 499.310 556.305 499.610 ;
        RECT 555.030 499.300 555.410 499.310 ;
        RECT 555.975 499.295 556.305 499.310 ;
        RECT 552.065 482.610 552.395 482.625 ;
        RECT 555.030 482.610 555.410 482.620 ;
        RECT 552.065 482.310 555.410 482.610 ;
        RECT 552.065 482.295 552.395 482.310 ;
        RECT 555.030 482.300 555.410 482.310 ;
      LAYER via3 ;
        RECT 555.060 499.300 555.380 499.620 ;
        RECT 555.060 482.300 555.380 482.620 ;
      LAYER met4 ;
        RECT 555.055 499.295 555.385 499.625 ;
        RECT 555.070 482.625 555.370 499.295 ;
        RECT 555.055 482.295 555.385 482.625 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 404.870 750.960 405.190 751.020 ;
        RECT 457.540 750.960 457.860 751.020 ;
        RECT 404.870 750.820 457.860 750.960 ;
        RECT 404.870 750.760 405.190 750.820 ;
        RECT 457.540 750.760 457.860 750.820 ;
        RECT 404.870 481.680 405.190 481.740 ;
        RECT 468.810 481.680 469.130 481.740 ;
        RECT 472.950 481.680 473.270 481.740 ;
        RECT 404.870 481.540 473.270 481.680 ;
        RECT 404.870 481.480 405.190 481.540 ;
        RECT 468.810 481.480 469.130 481.540 ;
        RECT 472.950 481.480 473.270 481.540 ;
        RECT 472.950 453.460 473.270 453.520 ;
        RECT 793.570 453.460 793.890 453.520 ;
        RECT 472.950 453.320 793.890 453.460 ;
        RECT 472.950 453.260 473.270 453.320 ;
        RECT 793.570 453.260 793.890 453.320 ;
      LAYER via ;
        RECT 404.900 750.760 405.160 751.020 ;
        RECT 457.570 750.760 457.830 751.020 ;
        RECT 404.900 481.480 405.160 481.740 ;
        RECT 468.840 481.480 469.100 481.740 ;
        RECT 472.980 481.480 473.240 481.740 ;
        RECT 472.980 453.260 473.240 453.520 ;
        RECT 793.600 453.260 793.860 453.520 ;
      LAYER met2 ;
        RECT 404.900 750.730 405.160 751.050 ;
        RECT 457.570 750.730 457.830 751.050 ;
        RECT 404.960 481.770 405.100 750.730 ;
        RECT 457.630 750.000 457.770 750.730 ;
        RECT 457.590 746.000 457.870 750.000 ;
        RECT 469.090 500.000 469.370 504.000 ;
        RECT 469.130 499.700 469.270 500.000 ;
        RECT 468.900 499.560 469.270 499.700 ;
        RECT 468.900 481.770 469.040 499.560 ;
        RECT 404.900 481.450 405.160 481.770 ;
        RECT 468.840 481.450 469.100 481.770 ;
        RECT 472.980 481.450 473.240 481.770 ;
        RECT 473.040 453.550 473.180 481.450 ;
        RECT 472.980 453.230 473.240 453.550 ;
        RECT 793.600 453.230 793.860 453.550 ;
        RECT 793.660 17.410 793.800 453.230 ;
        RECT 793.660 17.270 794.720 17.410 ;
        RECT 794.580 2.400 794.720 17.270 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 557.360 499.160 557.680 499.420 ;
        RECT 557.450 498.740 557.590 499.160 ;
        RECT 557.130 498.540 557.590 498.740 ;
        RECT 557.130 498.480 557.450 498.540 ;
      LAYER via ;
        RECT 557.390 499.160 557.650 499.420 ;
        RECT 557.160 498.480 557.420 498.740 ;
      LAYER met2 ;
        RECT 557.410 500.000 557.690 504.000 ;
        RECT 557.450 499.450 557.590 500.000 ;
        RECT 557.390 499.130 557.650 499.450 ;
        RECT 557.160 498.450 557.420 498.770 ;
        RECT 557.220 477.885 557.360 498.450 ;
        RECT 557.150 477.515 557.430 477.885 ;
        RECT 1854.350 74.275 1854.630 74.645 ;
        RECT 1854.420 2.400 1854.560 74.275 ;
        RECT 1854.210 -4.800 1854.770 2.400 ;
      LAYER via2 ;
        RECT 557.150 477.560 557.430 477.840 ;
        RECT 1854.350 74.320 1854.630 74.600 ;
      LAYER met3 ;
        RECT 557.125 477.860 557.455 477.865 ;
        RECT 556.870 477.850 557.455 477.860 ;
        RECT 556.670 477.550 557.455 477.850 ;
        RECT 556.870 477.540 557.455 477.550 ;
        RECT 557.125 477.535 557.455 477.540 ;
        RECT 556.870 74.610 557.250 74.620 ;
        RECT 1854.325 74.610 1854.655 74.625 ;
        RECT 556.870 74.310 1854.655 74.610 ;
        RECT 556.870 74.300 557.250 74.310 ;
        RECT 1854.325 74.295 1854.655 74.310 ;
      LAYER via3 ;
        RECT 556.900 477.540 557.220 477.860 ;
        RECT 556.900 74.300 557.220 74.620 ;
      LAYER met4 ;
        RECT 556.895 477.535 557.225 477.865 ;
        RECT 556.910 74.625 557.210 477.535 ;
        RECT 556.895 74.295 557.225 74.625 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.510 470.800 558.830 470.860 ;
        RECT 562.190 470.800 562.510 470.860 ;
        RECT 558.510 470.660 562.510 470.800 ;
        RECT 558.510 470.600 558.830 470.660 ;
        RECT 562.190 470.600 562.510 470.660 ;
        RECT 562.190 198.120 562.510 198.180 ;
        RECT 1870.430 198.120 1870.750 198.180 ;
        RECT 562.190 197.980 1870.750 198.120 ;
        RECT 562.190 197.920 562.510 197.980 ;
        RECT 1870.430 197.920 1870.750 197.980 ;
      LAYER via ;
        RECT 558.540 470.600 558.800 470.860 ;
        RECT 562.220 470.600 562.480 470.860 ;
        RECT 562.220 197.920 562.480 198.180 ;
        RECT 1870.460 197.920 1870.720 198.180 ;
      LAYER met2 ;
        RECT 558.790 500.000 559.070 504.000 ;
        RECT 558.830 499.645 558.970 500.000 ;
        RECT 558.760 499.275 559.040 499.645 ;
        RECT 558.530 498.850 558.810 498.965 ;
        RECT 558.530 498.710 559.200 498.850 ;
        RECT 558.530 498.595 558.810 498.710 ;
        RECT 559.060 473.690 559.200 498.710 ;
        RECT 558.600 473.550 559.200 473.690 ;
        RECT 558.600 470.890 558.740 473.550 ;
        RECT 558.540 470.570 558.800 470.890 ;
        RECT 562.220 470.570 562.480 470.890 ;
        RECT 562.280 198.210 562.420 470.570 ;
        RECT 562.220 197.890 562.480 198.210 ;
        RECT 1870.460 197.890 1870.720 198.210 ;
        RECT 1870.520 82.870 1870.660 197.890 ;
        RECT 1870.520 82.730 1871.120 82.870 ;
        RECT 1870.980 2.400 1871.120 82.730 ;
        RECT 1870.770 -4.800 1871.330 2.400 ;
      LAYER via2 ;
        RECT 558.760 499.320 559.040 499.600 ;
        RECT 558.530 498.640 558.810 498.920 ;
      LAYER met3 ;
        RECT 558.735 499.295 559.065 499.625 ;
        RECT 558.750 498.945 559.050 499.295 ;
        RECT 558.505 498.630 559.050 498.945 ;
        RECT 558.505 498.615 558.835 498.630 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.120 499.500 560.440 499.760 ;
        RECT 560.210 498.400 560.350 499.500 ;
        RECT 559.890 498.200 560.350 498.400 ;
        RECT 559.890 498.140 560.210 498.200 ;
        RECT 560.350 472.840 560.670 472.900 ;
        RECT 560.350 472.700 563.340 472.840 ;
        RECT 560.350 472.640 560.670 472.700 ;
        RECT 562.650 471.140 562.970 471.200 ;
        RECT 563.200 471.140 563.340 472.700 ;
        RECT 562.650 471.000 563.340 471.140 ;
        RECT 562.650 470.940 562.970 471.000 ;
        RECT 562.650 425.240 562.970 425.300 ;
        RECT 1883.770 425.240 1884.090 425.300 ;
        RECT 562.650 425.100 1884.090 425.240 ;
        RECT 562.650 425.040 562.970 425.100 ;
        RECT 1883.770 425.040 1884.090 425.100 ;
      LAYER via ;
        RECT 560.150 499.500 560.410 499.760 ;
        RECT 559.920 498.140 560.180 498.400 ;
        RECT 560.380 472.640 560.640 472.900 ;
        RECT 562.680 470.940 562.940 471.200 ;
        RECT 562.680 425.040 562.940 425.300 ;
        RECT 1883.800 425.040 1884.060 425.300 ;
      LAYER met2 ;
        RECT 560.170 500.000 560.450 504.000 ;
        RECT 560.210 499.790 560.350 500.000 ;
        RECT 560.150 499.470 560.410 499.790 ;
        RECT 559.920 498.110 560.180 498.430 ;
        RECT 559.980 497.490 560.120 498.110 ;
        RECT 559.980 497.350 560.580 497.490 ;
        RECT 560.440 472.930 560.580 497.350 ;
        RECT 560.380 472.610 560.640 472.930 ;
        RECT 562.680 470.910 562.940 471.230 ;
        RECT 562.740 425.330 562.880 470.910 ;
        RECT 562.680 425.010 562.940 425.330 ;
        RECT 1883.800 425.010 1884.060 425.330 ;
        RECT 1883.860 82.870 1884.000 425.010 ;
        RECT 1883.860 82.730 1887.680 82.870 ;
        RECT 1887.540 2.400 1887.680 82.730 ;
        RECT 1887.330 -4.800 1887.890 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.500 499.160 561.820 499.420 ;
        RECT 561.590 496.980 561.730 499.160 ;
        RECT 563.110 496.980 563.430 497.040 ;
        RECT 561.590 496.840 563.430 496.980 ;
        RECT 563.110 496.780 563.430 496.840 ;
        RECT 563.110 424.900 563.430 424.960 ;
        RECT 1897.570 424.900 1897.890 424.960 ;
        RECT 563.110 424.760 1897.890 424.900 ;
        RECT 563.110 424.700 563.430 424.760 ;
        RECT 1897.570 424.700 1897.890 424.760 ;
        RECT 1897.570 16.900 1897.890 16.960 ;
        RECT 1904.010 16.900 1904.330 16.960 ;
        RECT 1897.570 16.760 1904.330 16.900 ;
        RECT 1897.570 16.700 1897.890 16.760 ;
        RECT 1904.010 16.700 1904.330 16.760 ;
      LAYER via ;
        RECT 561.530 499.160 561.790 499.420 ;
        RECT 563.140 496.780 563.400 497.040 ;
        RECT 563.140 424.700 563.400 424.960 ;
        RECT 1897.600 424.700 1897.860 424.960 ;
        RECT 1897.600 16.700 1897.860 16.960 ;
        RECT 1904.040 16.700 1904.300 16.960 ;
      LAYER met2 ;
        RECT 561.550 500.000 561.830 504.000 ;
        RECT 561.590 499.450 561.730 500.000 ;
        RECT 561.530 499.130 561.790 499.450 ;
        RECT 563.140 496.750 563.400 497.070 ;
        RECT 563.200 424.990 563.340 496.750 ;
        RECT 563.140 424.670 563.400 424.990 ;
        RECT 1897.600 424.670 1897.860 424.990 ;
        RECT 1897.660 16.990 1897.800 424.670 ;
        RECT 1897.600 16.670 1897.860 16.990 ;
        RECT 1904.040 16.670 1904.300 16.990 ;
        RECT 1904.100 2.400 1904.240 16.670 ;
        RECT 1903.890 -4.800 1904.450 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.880 500.180 563.200 500.440 ;
        RECT 562.970 499.700 563.110 500.180 ;
        RECT 561.130 499.560 563.110 499.700 ;
        RECT 559.890 496.980 560.210 497.040 ;
        RECT 561.130 496.980 561.270 499.560 ;
        RECT 559.890 496.840 561.270 496.980 ;
        RECT 559.890 496.780 560.210 496.840 ;
        RECT 558.970 472.840 559.290 472.900 ;
        RECT 559.890 472.840 560.210 472.900 ;
        RECT 558.970 472.700 560.210 472.840 ;
        RECT 558.970 472.640 559.290 472.700 ;
        RECT 559.890 472.640 560.210 472.700 ;
        RECT 558.970 73.340 559.290 73.400 ;
        RECT 1920.570 73.340 1920.890 73.400 ;
        RECT 558.970 73.200 1920.890 73.340 ;
        RECT 558.970 73.140 559.290 73.200 ;
        RECT 1920.570 73.140 1920.890 73.200 ;
      LAYER via ;
        RECT 562.910 500.180 563.170 500.440 ;
        RECT 559.920 496.780 560.180 497.040 ;
        RECT 559.000 472.640 559.260 472.900 ;
        RECT 559.920 472.640 560.180 472.900 ;
        RECT 559.000 73.140 559.260 73.400 ;
        RECT 1920.600 73.140 1920.860 73.400 ;
      LAYER met2 ;
        RECT 562.930 500.470 563.210 504.000 ;
        RECT 562.910 500.150 563.210 500.470 ;
        RECT 562.930 500.000 563.210 500.150 ;
        RECT 559.920 496.750 560.180 497.070 ;
        RECT 559.980 472.930 560.120 496.750 ;
        RECT 559.000 472.610 559.260 472.930 ;
        RECT 559.920 472.610 560.180 472.930 ;
        RECT 559.060 73.430 559.200 472.610 ;
        RECT 559.000 73.110 559.260 73.430 ;
        RECT 1920.600 73.110 1920.860 73.430 ;
        RECT 1920.660 2.400 1920.800 73.110 ;
        RECT 1920.450 -4.800 1921.010 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.310 500.000 564.590 504.000 ;
        RECT 564.350 498.340 564.490 500.000 ;
        RECT 564.120 498.200 564.490 498.340 ;
        RECT 564.120 484.685 564.260 498.200 ;
        RECT 564.050 484.315 564.330 484.685 ;
        RECT 1937.150 72.915 1937.430 73.285 ;
        RECT 1937.220 2.400 1937.360 72.915 ;
        RECT 1937.010 -4.800 1937.570 2.400 ;
      LAYER via2 ;
        RECT 564.050 484.360 564.330 484.640 ;
        RECT 1937.150 72.960 1937.430 73.240 ;
      LAYER met3 ;
        RECT 564.025 484.650 564.355 484.665 ;
        RECT 565.150 484.650 565.530 484.660 ;
        RECT 564.025 484.350 565.530 484.650 ;
        RECT 564.025 484.335 564.355 484.350 ;
        RECT 565.150 484.340 565.530 484.350 ;
        RECT 565.150 73.250 565.530 73.260 ;
        RECT 1937.125 73.250 1937.455 73.265 ;
        RECT 565.150 72.950 1937.455 73.250 ;
        RECT 565.150 72.940 565.530 72.950 ;
        RECT 1937.125 72.935 1937.455 72.950 ;
      LAYER via3 ;
        RECT 565.180 484.340 565.500 484.660 ;
        RECT 565.180 72.940 565.500 73.260 ;
      LAYER met4 ;
        RECT 565.175 484.335 565.505 484.665 ;
        RECT 565.190 73.265 565.490 484.335 ;
        RECT 565.175 72.935 565.505 73.265 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.640 499.160 565.960 499.420 ;
        RECT 565.730 498.000 565.870 499.160 ;
        RECT 567.250 498.000 567.570 498.060 ;
        RECT 565.730 497.860 567.570 498.000 ;
        RECT 567.250 497.800 567.570 497.860 ;
        RECT 567.250 475.220 567.570 475.280 ;
        RECT 569.090 475.220 569.410 475.280 ;
        RECT 567.250 475.080 569.410 475.220 ;
        RECT 567.250 475.020 567.570 475.080 ;
        RECT 569.090 475.020 569.410 475.080 ;
        RECT 569.090 410.960 569.410 411.020 ;
        RECT 1952.770 410.960 1953.090 411.020 ;
        RECT 569.090 410.820 1953.090 410.960 ;
        RECT 569.090 410.760 569.410 410.820 ;
        RECT 1952.770 410.760 1953.090 410.820 ;
      LAYER via ;
        RECT 565.670 499.160 565.930 499.420 ;
        RECT 567.280 497.800 567.540 498.060 ;
        RECT 567.280 475.020 567.540 475.280 ;
        RECT 569.120 475.020 569.380 475.280 ;
        RECT 569.120 410.760 569.380 411.020 ;
        RECT 1952.800 410.760 1953.060 411.020 ;
      LAYER met2 ;
        RECT 565.690 500.000 565.970 504.000 ;
        RECT 565.730 499.450 565.870 500.000 ;
        RECT 565.670 499.130 565.930 499.450 ;
        RECT 567.280 497.770 567.540 498.090 ;
        RECT 567.340 475.310 567.480 497.770 ;
        RECT 567.280 474.990 567.540 475.310 ;
        RECT 569.120 474.990 569.380 475.310 ;
        RECT 569.180 411.050 569.320 474.990 ;
        RECT 569.120 410.730 569.380 411.050 ;
        RECT 1952.800 410.730 1953.060 411.050 ;
        RECT 1952.860 17.410 1953.000 410.730 ;
        RECT 1952.860 17.270 1953.920 17.410 ;
        RECT 1953.780 2.400 1953.920 17.270 ;
        RECT 1953.570 -4.800 1954.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 73.000 567.110 73.060 ;
        RECT 1970.250 73.000 1970.570 73.060 ;
        RECT 566.790 72.860 1970.570 73.000 ;
        RECT 566.790 72.800 567.110 72.860 ;
        RECT 1970.250 72.800 1970.570 72.860 ;
      LAYER via ;
        RECT 566.820 72.800 567.080 73.060 ;
        RECT 1970.280 72.800 1970.540 73.060 ;
      LAYER met2 ;
        RECT 567.070 500.000 567.350 504.000 ;
        RECT 567.110 498.850 567.250 500.000 ;
        RECT 566.880 498.710 567.250 498.850 ;
        RECT 566.880 73.090 567.020 498.710 ;
        RECT 566.820 72.770 567.080 73.090 ;
        RECT 1970.280 72.770 1970.540 73.090 ;
        RECT 1970.340 2.400 1970.480 72.770 ;
        RECT 1970.130 -4.800 1970.690 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.400 499.700 568.720 499.760 ;
        RECT 567.110 499.560 568.720 499.700 ;
        RECT 566.330 498.340 566.650 498.400 ;
        RECT 567.110 498.340 567.250 499.560 ;
        RECT 568.400 499.500 568.720 499.560 ;
        RECT 566.330 498.200 567.250 498.340 ;
        RECT 566.330 498.140 566.650 498.200 ;
        RECT 565.870 72.660 566.190 72.720 ;
        RECT 1980.830 72.660 1981.150 72.720 ;
        RECT 565.870 72.520 1981.150 72.660 ;
        RECT 565.870 72.460 566.190 72.520 ;
        RECT 1980.830 72.460 1981.150 72.520 ;
        RECT 1980.830 20.300 1981.150 20.360 ;
        RECT 1986.810 20.300 1987.130 20.360 ;
        RECT 1980.830 20.160 1987.130 20.300 ;
        RECT 1980.830 20.100 1981.150 20.160 ;
        RECT 1986.810 20.100 1987.130 20.160 ;
      LAYER via ;
        RECT 566.360 498.140 566.620 498.400 ;
        RECT 568.430 499.500 568.690 499.760 ;
        RECT 565.900 72.460 566.160 72.720 ;
        RECT 1980.860 72.460 1981.120 72.720 ;
        RECT 1980.860 20.100 1981.120 20.360 ;
        RECT 1986.840 20.100 1987.100 20.360 ;
      LAYER met2 ;
        RECT 568.450 500.000 568.730 504.000 ;
        RECT 568.490 499.790 568.630 500.000 ;
        RECT 568.430 499.470 568.690 499.790 ;
        RECT 566.360 498.110 566.620 498.430 ;
        RECT 566.420 473.010 566.560 498.110 ;
        RECT 565.960 472.870 566.560 473.010 ;
        RECT 565.960 72.750 566.100 472.870 ;
        RECT 565.900 72.430 566.160 72.750 ;
        RECT 1980.860 72.430 1981.120 72.750 ;
        RECT 1980.920 20.390 1981.060 72.430 ;
        RECT 1980.860 20.070 1981.120 20.390 ;
        RECT 1986.840 20.070 1987.100 20.390 ;
        RECT 1986.900 2.400 1987.040 20.070 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 569.550 498.340 569.870 498.400 ;
        RECT 570.470 498.340 570.790 498.400 ;
        RECT 569.550 498.200 570.790 498.340 ;
        RECT 569.550 498.140 569.870 498.200 ;
        RECT 570.470 498.140 570.790 498.200 ;
        RECT 566.330 472.160 566.650 472.220 ;
        RECT 570.470 472.160 570.790 472.220 ;
        RECT 566.330 472.020 570.790 472.160 ;
        RECT 566.330 471.960 566.650 472.020 ;
        RECT 570.470 471.960 570.790 472.020 ;
        RECT 566.330 72.320 566.650 72.380 ;
        RECT 2003.370 72.320 2003.690 72.380 ;
        RECT 566.330 72.180 2003.690 72.320 ;
        RECT 566.330 72.120 566.650 72.180 ;
        RECT 2003.370 72.120 2003.690 72.180 ;
      LAYER via ;
        RECT 569.580 498.140 569.840 498.400 ;
        RECT 570.500 498.140 570.760 498.400 ;
        RECT 566.360 471.960 566.620 472.220 ;
        RECT 570.500 471.960 570.760 472.220 ;
        RECT 566.360 72.120 566.620 72.380 ;
        RECT 2003.400 72.120 2003.660 72.380 ;
      LAYER met2 ;
        RECT 569.830 500.000 570.110 504.000 ;
        RECT 569.870 499.530 570.010 500.000 ;
        RECT 569.640 499.390 570.010 499.530 ;
        RECT 569.640 498.430 569.780 499.390 ;
        RECT 569.580 498.110 569.840 498.430 ;
        RECT 570.500 498.110 570.760 498.430 ;
        RECT 570.560 472.250 570.700 498.110 ;
        RECT 566.360 471.930 566.620 472.250 ;
        RECT 570.500 471.930 570.760 472.250 ;
        RECT 566.420 72.410 566.560 471.930 ;
        RECT 566.360 72.090 566.620 72.410 ;
        RECT 2003.400 72.090 2003.660 72.410 ;
        RECT 2003.460 2.400 2003.600 72.090 ;
        RECT 2003.250 -4.800 2003.810 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 405.330 748.920 405.650 748.980 ;
        RECT 405.330 748.780 446.500 748.920 ;
        RECT 405.330 748.720 405.650 748.780 ;
        RECT 446.360 748.580 446.500 748.780 ;
        RECT 462.370 748.580 462.690 748.640 ;
        RECT 446.360 748.440 462.690 748.580 ;
        RECT 462.370 748.380 462.690 748.440 ;
        RECT 405.330 478.960 405.650 479.020 ;
        RECT 467.890 478.960 468.210 479.020 ;
        RECT 472.490 478.960 472.810 479.020 ;
        RECT 405.330 478.820 472.810 478.960 ;
        RECT 405.330 478.760 405.650 478.820 ;
        RECT 467.890 478.760 468.210 478.820 ;
        RECT 472.490 478.760 472.810 478.820 ;
        RECT 472.950 81.500 473.270 81.560 ;
        RECT 810.130 81.500 810.450 81.560 ;
        RECT 472.950 81.360 810.450 81.500 ;
        RECT 472.950 81.300 473.270 81.360 ;
        RECT 810.130 81.300 810.450 81.360 ;
      LAYER via ;
        RECT 405.360 748.720 405.620 748.980 ;
        RECT 462.400 748.380 462.660 748.640 ;
        RECT 405.360 478.760 405.620 479.020 ;
        RECT 467.920 478.760 468.180 479.020 ;
        RECT 472.520 478.760 472.780 479.020 ;
        RECT 472.980 81.300 473.240 81.560 ;
        RECT 810.160 81.300 810.420 81.560 ;
      LAYER met2 ;
        RECT 405.360 748.690 405.620 749.010 ;
        RECT 405.420 479.050 405.560 748.690 ;
        RECT 462.400 748.410 462.660 748.670 ;
        RECT 463.110 748.410 463.390 750.000 ;
        RECT 462.400 748.350 463.390 748.410 ;
        RECT 462.460 748.270 463.390 748.350 ;
        RECT 463.110 746.000 463.390 748.270 ;
        RECT 470.470 500.000 470.750 504.000 ;
        RECT 470.510 498.680 470.650 500.000 ;
        RECT 470.280 498.540 470.650 498.680 ;
        RECT 470.280 498.285 470.420 498.540 ;
        RECT 468.370 497.915 468.650 498.285 ;
        RECT 470.210 497.915 470.490 498.285 ;
        RECT 468.440 487.970 468.580 497.915 ;
        RECT 467.980 487.830 468.580 487.970 ;
        RECT 467.980 479.050 468.120 487.830 ;
        RECT 405.360 478.730 405.620 479.050 ;
        RECT 467.920 478.730 468.180 479.050 ;
        RECT 472.520 478.730 472.780 479.050 ;
        RECT 472.580 448.570 472.720 478.730 ;
        RECT 472.580 448.430 473.180 448.570 ;
        RECT 473.040 81.590 473.180 448.430 ;
        RECT 472.980 81.270 473.240 81.590 ;
        RECT 810.160 81.270 810.420 81.590 ;
        RECT 810.220 17.410 810.360 81.270 ;
        RECT 810.220 17.270 811.280 17.410 ;
        RECT 811.140 2.400 811.280 17.270 ;
        RECT 810.930 -4.800 811.490 2.400 ;
      LAYER via2 ;
        RECT 468.370 497.960 468.650 498.240 ;
        RECT 470.210 497.960 470.490 498.240 ;
      LAYER met3 ;
        RECT 468.345 498.250 468.675 498.265 ;
        RECT 470.185 498.250 470.515 498.265 ;
        RECT 468.345 497.950 470.515 498.250 ;
        RECT 468.345 497.935 468.675 497.950 ;
        RECT 470.185 497.935 470.515 497.950 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.210 500.000 571.490 504.000 ;
        RECT 571.250 498.850 571.390 500.000 ;
        RECT 571.020 498.710 571.390 498.850 ;
        RECT 571.020 484.005 571.160 498.710 ;
        RECT 570.950 483.635 571.230 484.005 ;
        RECT 2019.950 80.395 2020.230 80.765 ;
        RECT 2020.020 2.400 2020.160 80.395 ;
        RECT 2019.810 -4.800 2020.370 2.400 ;
      LAYER via2 ;
        RECT 570.950 483.680 571.230 483.960 ;
        RECT 2019.950 80.440 2020.230 80.720 ;
      LAYER met3 ;
        RECT 569.750 483.970 570.130 483.980 ;
        RECT 570.925 483.970 571.255 483.985 ;
        RECT 569.750 483.670 571.255 483.970 ;
        RECT 569.750 483.660 570.130 483.670 ;
        RECT 570.925 483.655 571.255 483.670 ;
        RECT 569.750 80.730 570.130 80.740 ;
        RECT 2019.925 80.730 2020.255 80.745 ;
        RECT 569.750 80.430 2020.255 80.730 ;
        RECT 569.750 80.420 570.130 80.430 ;
        RECT 2019.925 80.415 2020.255 80.430 ;
      LAYER via3 ;
        RECT 569.780 483.660 570.100 483.980 ;
        RECT 569.780 80.420 570.100 80.740 ;
      LAYER met4 ;
        RECT 569.775 483.655 570.105 483.985 ;
        RECT 569.790 80.745 570.090 483.655 ;
        RECT 569.775 80.415 570.105 80.745 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.450 439.860 576.770 439.920 ;
        RECT 2035.570 439.860 2035.890 439.920 ;
        RECT 576.450 439.720 2035.890 439.860 ;
        RECT 576.450 439.660 576.770 439.720 ;
        RECT 2035.570 439.660 2035.890 439.720 ;
      LAYER via ;
        RECT 576.480 439.660 576.740 439.920 ;
        RECT 2035.600 439.660 2035.860 439.920 ;
      LAYER met2 ;
        RECT 572.590 500.000 572.870 504.000 ;
        RECT 572.630 499.645 572.770 500.000 ;
        RECT 572.560 499.275 572.840 499.645 ;
        RECT 576.010 496.615 576.290 496.985 ;
        RECT 576.080 473.010 576.220 496.615 ;
        RECT 576.080 472.870 576.680 473.010 ;
        RECT 576.540 439.950 576.680 472.870 ;
        RECT 576.480 439.630 576.740 439.950 ;
        RECT 2035.600 439.630 2035.860 439.950 ;
        RECT 2035.660 17.410 2035.800 439.630 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
      LAYER via2 ;
        RECT 572.560 499.320 572.840 499.600 ;
        RECT 576.010 496.660 576.290 496.940 ;
      LAYER met3 ;
        RECT 572.535 499.610 572.865 499.625 ;
        RECT 572.535 499.310 576.530 499.610 ;
        RECT 572.535 499.295 572.865 499.310 ;
        RECT 576.230 496.965 576.530 499.310 ;
        RECT 575.985 496.650 576.530 496.965 ;
        RECT 575.985 496.635 576.315 496.650 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 475.900 574.470 475.960 ;
        RECT 577.370 475.900 577.690 475.960 ;
        RECT 574.150 475.760 577.690 475.900 ;
        RECT 574.150 475.700 574.470 475.760 ;
        RECT 577.370 475.700 577.690 475.760 ;
        RECT 576.910 445.300 577.230 445.360 ;
        RECT 2049.370 445.300 2049.690 445.360 ;
        RECT 576.910 445.160 2049.690 445.300 ;
        RECT 576.910 445.100 577.230 445.160 ;
        RECT 2049.370 445.100 2049.690 445.160 ;
      LAYER via ;
        RECT 574.180 475.700 574.440 475.960 ;
        RECT 577.400 475.700 577.660 475.960 ;
        RECT 576.940 445.100 577.200 445.360 ;
        RECT 2049.400 445.100 2049.660 445.360 ;
      LAYER met2 ;
        RECT 573.970 500.000 574.250 504.000 ;
        RECT 574.010 498.680 574.150 500.000 ;
        RECT 573.780 498.540 574.150 498.680 ;
        RECT 573.780 497.660 573.920 498.540 ;
        RECT 573.780 497.520 574.380 497.660 ;
        RECT 574.240 475.990 574.380 497.520 ;
        RECT 574.180 475.670 574.440 475.990 ;
        RECT 577.400 475.670 577.660 475.990 ;
        RECT 577.460 448.570 577.600 475.670 ;
        RECT 577.000 448.430 577.600 448.570 ;
        RECT 577.000 445.390 577.140 448.430 ;
        RECT 576.940 445.070 577.200 445.390 ;
        RECT 2049.400 445.070 2049.660 445.390 ;
        RECT 2049.460 82.870 2049.600 445.070 ;
        RECT 2049.460 82.730 2053.280 82.870 ;
        RECT 2053.140 2.400 2053.280 82.730 ;
        RECT 2052.930 -4.800 2053.490 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.230 81.160 573.550 81.220 ;
        RECT 2063.630 81.160 2063.950 81.220 ;
        RECT 573.230 81.020 2063.950 81.160 ;
        RECT 573.230 80.960 573.550 81.020 ;
        RECT 2063.630 80.960 2063.950 81.020 ;
        RECT 2063.630 16.900 2063.950 16.960 ;
        RECT 2069.610 16.900 2069.930 16.960 ;
        RECT 2063.630 16.760 2069.930 16.900 ;
        RECT 2063.630 16.700 2063.950 16.760 ;
        RECT 2069.610 16.700 2069.930 16.760 ;
      LAYER via ;
        RECT 573.260 80.960 573.520 81.220 ;
        RECT 2063.660 80.960 2063.920 81.220 ;
        RECT 2063.660 16.700 2063.920 16.960 ;
        RECT 2069.640 16.700 2069.900 16.960 ;
      LAYER met2 ;
        RECT 575.350 500.000 575.630 504.000 ;
        RECT 575.390 498.850 575.530 500.000 ;
        RECT 575.160 498.795 575.530 498.850 ;
        RECT 575.090 498.710 575.530 498.795 ;
        RECT 575.090 498.425 575.370 498.710 ;
        RECT 573.250 497.915 573.530 498.285 ;
        RECT 573.320 81.250 573.460 497.915 ;
        RECT 573.260 80.930 573.520 81.250 ;
        RECT 2063.660 80.930 2063.920 81.250 ;
        RECT 2063.720 16.990 2063.860 80.930 ;
        RECT 2063.660 16.670 2063.920 16.990 ;
        RECT 2069.640 16.670 2069.900 16.990 ;
        RECT 2069.700 2.400 2069.840 16.670 ;
        RECT 2069.490 -4.800 2070.050 2.400 ;
      LAYER via2 ;
        RECT 575.090 498.470 575.370 498.750 ;
        RECT 573.250 497.960 573.530 498.240 ;
      LAYER met3 ;
        RECT 573.470 498.630 575.610 498.930 ;
        RECT 573.470 498.265 573.770 498.630 ;
        RECT 575.065 498.460 575.610 498.630 ;
        RECT 575.065 498.445 575.395 498.460 ;
        RECT 573.225 497.950 573.770 498.265 ;
        RECT 573.225 497.935 573.555 497.950 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.680 499.500 577.000 499.760 ;
        RECT 576.770 497.720 576.910 499.500 ;
        RECT 576.770 497.520 577.230 497.720 ;
        RECT 576.910 497.460 577.230 497.520 ;
        RECT 573.690 471.820 574.010 471.880 ;
        RECT 577.830 471.820 578.150 471.880 ;
        RECT 573.690 471.680 578.150 471.820 ;
        RECT 573.690 471.620 574.010 471.680 ;
        RECT 577.830 471.620 578.150 471.680 ;
        RECT 573.690 80.820 574.010 80.880 ;
        RECT 2086.170 80.820 2086.490 80.880 ;
        RECT 573.690 80.680 2086.490 80.820 ;
        RECT 573.690 80.620 574.010 80.680 ;
        RECT 2086.170 80.620 2086.490 80.680 ;
      LAYER via ;
        RECT 576.710 499.500 576.970 499.760 ;
        RECT 576.940 497.460 577.200 497.720 ;
        RECT 573.720 471.620 573.980 471.880 ;
        RECT 577.860 471.620 578.120 471.880 ;
        RECT 573.720 80.620 573.980 80.880 ;
        RECT 2086.200 80.620 2086.460 80.880 ;
      LAYER met2 ;
        RECT 576.730 500.000 577.010 504.000 ;
        RECT 576.770 499.790 576.910 500.000 ;
        RECT 576.710 499.470 576.970 499.790 ;
        RECT 576.940 497.430 577.200 497.750 ;
        RECT 577.000 476.410 577.140 497.430 ;
        RECT 577.000 476.270 578.060 476.410 ;
        RECT 577.920 471.910 578.060 476.270 ;
        RECT 573.720 471.590 573.980 471.910 ;
        RECT 577.860 471.590 578.120 471.910 ;
        RECT 573.780 80.910 573.920 471.590 ;
        RECT 573.720 80.590 573.980 80.910 ;
        RECT 2086.200 80.590 2086.460 80.910 ;
        RECT 2086.260 2.400 2086.400 80.590 ;
        RECT 2086.050 -4.800 2086.610 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.110 500.000 578.390 504.000 ;
        RECT 578.150 498.340 578.290 500.000 ;
        RECT 577.920 498.200 578.290 498.340 ;
        RECT 577.920 483.325 578.060 498.200 ;
        RECT 577.850 482.955 578.130 483.325 ;
        RECT 2102.750 79.035 2103.030 79.405 ;
        RECT 2102.820 2.400 2102.960 79.035 ;
        RECT 2102.610 -4.800 2103.170 2.400 ;
      LAYER via2 ;
        RECT 577.850 483.000 578.130 483.280 ;
        RECT 2102.750 79.080 2103.030 79.360 ;
      LAYER met3 ;
        RECT 577.825 483.290 578.155 483.305 ;
        RECT 578.950 483.290 579.330 483.300 ;
        RECT 577.825 482.990 579.330 483.290 ;
        RECT 577.825 482.975 578.155 482.990 ;
        RECT 578.950 482.980 579.330 482.990 ;
        RECT 578.950 79.370 579.330 79.380 ;
        RECT 2102.725 79.370 2103.055 79.385 ;
        RECT 578.950 79.070 2103.055 79.370 ;
        RECT 578.950 79.060 579.330 79.070 ;
        RECT 2102.725 79.055 2103.055 79.070 ;
      LAYER via3 ;
        RECT 578.980 482.980 579.300 483.300 ;
        RECT 578.980 79.060 579.300 79.380 ;
      LAYER met4 ;
        RECT 578.975 482.975 579.305 483.305 ;
        RECT 578.990 79.385 579.290 482.975 ;
        RECT 578.975 79.055 579.305 79.385 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.440 499.500 579.760 499.760 ;
        RECT 579.530 498.000 579.670 499.500 ;
        RECT 580.130 498.000 580.450 498.060 ;
        RECT 579.530 497.860 580.450 498.000 ;
        RECT 580.130 497.800 580.450 497.860 ;
        RECT 580.130 475.220 580.450 475.280 ;
        RECT 581.970 475.220 582.290 475.280 ;
        RECT 580.130 475.080 582.290 475.220 ;
        RECT 580.130 475.020 580.450 475.080 ;
        RECT 581.970 475.020 582.290 475.080 ;
        RECT 581.970 204.580 582.290 204.640 ;
        RECT 2118.370 204.580 2118.690 204.640 ;
        RECT 581.970 204.440 2118.690 204.580 ;
        RECT 581.970 204.380 582.290 204.440 ;
        RECT 2118.370 204.380 2118.690 204.440 ;
      LAYER via ;
        RECT 579.470 499.500 579.730 499.760 ;
        RECT 580.160 497.800 580.420 498.060 ;
        RECT 580.160 475.020 580.420 475.280 ;
        RECT 582.000 475.020 582.260 475.280 ;
        RECT 582.000 204.380 582.260 204.640 ;
        RECT 2118.400 204.380 2118.660 204.640 ;
      LAYER met2 ;
        RECT 579.490 500.000 579.770 504.000 ;
        RECT 579.530 499.790 579.670 500.000 ;
        RECT 579.470 499.470 579.730 499.790 ;
        RECT 580.160 497.770 580.420 498.090 ;
        RECT 580.220 475.310 580.360 497.770 ;
        RECT 580.160 474.990 580.420 475.310 ;
        RECT 582.000 474.990 582.260 475.310 ;
        RECT 582.060 204.670 582.200 474.990 ;
        RECT 582.000 204.350 582.260 204.670 ;
        RECT 2118.400 204.350 2118.660 204.670 ;
        RECT 2118.460 17.410 2118.600 204.350 ;
        RECT 2118.460 17.270 2119.520 17.410 ;
        RECT 2119.380 2.400 2119.520 17.270 ;
        RECT 2119.170 -4.800 2119.730 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.430 424.560 582.750 424.620 ;
        RECT 2132.170 424.560 2132.490 424.620 ;
        RECT 582.430 424.420 2132.490 424.560 ;
        RECT 582.430 424.360 582.750 424.420 ;
        RECT 2132.170 424.360 2132.490 424.420 ;
      LAYER via ;
        RECT 582.460 424.360 582.720 424.620 ;
        RECT 2132.200 424.360 2132.460 424.620 ;
      LAYER met2 ;
        RECT 580.870 500.000 581.150 504.000 ;
        RECT 580.910 499.815 581.050 500.000 ;
        RECT 580.840 499.445 581.120 499.815 ;
        RECT 581.990 498.595 582.270 498.965 ;
        RECT 582.060 487.970 582.200 498.595 ;
        RECT 582.060 487.830 582.660 487.970 ;
        RECT 582.520 424.650 582.660 487.830 ;
        RECT 582.460 424.330 582.720 424.650 ;
        RECT 2132.200 424.330 2132.460 424.650 ;
        RECT 2132.260 82.870 2132.400 424.330 ;
        RECT 2132.260 82.730 2136.080 82.870 ;
        RECT 2135.940 2.400 2136.080 82.730 ;
        RECT 2135.730 -4.800 2136.290 2.400 ;
      LAYER via2 ;
        RECT 580.840 499.490 581.120 499.770 ;
        RECT 581.990 498.640 582.270 498.920 ;
      LAYER met3 ;
        RECT 580.815 499.465 581.145 499.795 ;
        RECT 580.830 498.930 581.130 499.465 ;
        RECT 581.965 498.930 582.295 498.945 ;
        RECT 580.830 498.630 582.295 498.930 ;
        RECT 581.965 498.615 582.295 498.630 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 582.200 499.500 582.520 499.760 ;
        RECT 582.290 499.080 582.430 499.500 ;
        RECT 582.290 498.880 582.750 499.080 ;
        RECT 582.430 498.820 582.750 498.880 ;
        RECT 582.430 496.440 582.750 496.700 ;
        RECT 582.520 495.620 582.660 496.440 ;
        RECT 583.350 495.620 583.670 495.680 ;
        RECT 582.520 495.480 583.670 495.620 ;
        RECT 583.350 495.420 583.670 495.480 ;
        RECT 583.350 444.960 583.670 445.020 ;
        RECT 2145.970 444.960 2146.290 445.020 ;
        RECT 583.350 444.820 2146.290 444.960 ;
        RECT 583.350 444.760 583.670 444.820 ;
        RECT 2145.970 444.760 2146.290 444.820 ;
        RECT 2145.970 16.900 2146.290 16.960 ;
        RECT 2152.410 16.900 2152.730 16.960 ;
        RECT 2145.970 16.760 2152.730 16.900 ;
        RECT 2145.970 16.700 2146.290 16.760 ;
        RECT 2152.410 16.700 2152.730 16.760 ;
      LAYER via ;
        RECT 582.230 499.500 582.490 499.760 ;
        RECT 582.460 498.820 582.720 499.080 ;
        RECT 582.460 496.440 582.720 496.700 ;
        RECT 583.380 495.420 583.640 495.680 ;
        RECT 583.380 444.760 583.640 445.020 ;
        RECT 2146.000 444.760 2146.260 445.020 ;
        RECT 2146.000 16.700 2146.260 16.960 ;
        RECT 2152.440 16.700 2152.700 16.960 ;
      LAYER met2 ;
        RECT 582.250 500.000 582.530 504.000 ;
        RECT 582.290 499.790 582.430 500.000 ;
        RECT 582.230 499.470 582.490 499.790 ;
        RECT 582.460 498.790 582.720 499.110 ;
        RECT 582.520 496.730 582.660 498.790 ;
        RECT 582.460 496.410 582.720 496.730 ;
        RECT 583.380 495.390 583.640 495.710 ;
        RECT 583.440 445.050 583.580 495.390 ;
        RECT 583.380 444.730 583.640 445.050 ;
        RECT 2146.000 444.730 2146.260 445.050 ;
        RECT 2146.060 16.990 2146.200 444.730 ;
        RECT 2146.000 16.670 2146.260 16.990 ;
        RECT 2152.440 16.670 2152.700 16.990 ;
        RECT 2152.500 2.400 2152.640 16.670 ;
        RECT 2152.290 -4.800 2152.850 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.830 500.240 583.810 500.380 ;
        RECT 581.830 498.680 581.970 500.240 ;
        RECT 583.670 499.760 583.810 500.240 ;
        RECT 583.580 499.500 583.900 499.760 ;
        RECT 582.890 498.680 583.210 498.740 ;
        RECT 581.830 498.540 583.210 498.680 ;
        RECT 582.890 498.480 583.210 498.540 ;
        RECT 582.890 431.700 583.210 431.760 ;
        RECT 2166.670 431.700 2166.990 431.760 ;
        RECT 582.890 431.560 2166.990 431.700 ;
        RECT 582.890 431.500 583.210 431.560 ;
        RECT 2166.670 431.500 2166.990 431.560 ;
      LAYER via ;
        RECT 583.610 499.500 583.870 499.760 ;
        RECT 582.920 498.480 583.180 498.740 ;
        RECT 582.920 431.500 583.180 431.760 ;
        RECT 2166.700 431.500 2166.960 431.760 ;
      LAYER met2 ;
        RECT 583.630 500.000 583.910 504.000 ;
        RECT 583.670 499.790 583.810 500.000 ;
        RECT 583.610 499.470 583.870 499.790 ;
        RECT 582.920 498.450 583.180 498.770 ;
        RECT 582.980 431.790 583.120 498.450 ;
        RECT 582.920 431.470 583.180 431.790 ;
        RECT 2166.700 431.470 2166.960 431.790 ;
        RECT 2166.760 82.870 2166.900 431.470 ;
        RECT 2166.760 82.730 2169.200 82.870 ;
        RECT 2169.060 2.400 2169.200 82.730 ;
        RECT 2168.850 -4.800 2169.410 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 406.710 749.940 407.030 750.000 ;
        RECT 406.710 749.800 447.420 749.940 ;
        RECT 406.710 749.740 407.030 749.800 ;
        RECT 447.280 749.260 447.420 749.800 ;
        RECT 467.890 749.260 468.210 749.320 ;
        RECT 447.280 749.120 468.210 749.260 ;
        RECT 467.890 749.060 468.210 749.120 ;
        RECT 471.800 499.500 472.120 499.760 ;
        RECT 471.110 497.660 471.430 497.720 ;
        RECT 471.890 497.660 472.030 499.500 ;
        RECT 471.110 497.520 472.030 497.660 ;
        RECT 471.110 497.460 471.430 497.520 ;
        RECT 406.710 482.020 407.030 482.080 ;
        RECT 471.110 482.020 471.430 482.080 ;
        RECT 473.410 482.020 473.730 482.080 ;
        RECT 406.710 481.880 473.730 482.020 ;
        RECT 406.710 481.820 407.030 481.880 ;
        RECT 471.110 481.820 471.430 481.880 ;
        RECT 473.410 481.820 473.730 481.880 ;
        RECT 473.410 87.960 473.730 88.020 ;
        RECT 821.630 87.960 821.950 88.020 ;
        RECT 473.410 87.820 821.950 87.960 ;
        RECT 473.410 87.760 473.730 87.820 ;
        RECT 821.630 87.760 821.950 87.820 ;
        RECT 821.630 19.280 821.950 19.340 ;
        RECT 827.610 19.280 827.930 19.340 ;
        RECT 821.630 19.140 827.930 19.280 ;
        RECT 821.630 19.080 821.950 19.140 ;
        RECT 827.610 19.080 827.930 19.140 ;
      LAYER via ;
        RECT 406.740 749.740 407.000 750.000 ;
        RECT 467.920 749.060 468.180 749.320 ;
        RECT 471.830 499.500 472.090 499.760 ;
        RECT 471.140 497.460 471.400 497.720 ;
        RECT 406.740 481.820 407.000 482.080 ;
        RECT 471.140 481.820 471.400 482.080 ;
        RECT 473.440 481.820 473.700 482.080 ;
        RECT 473.440 87.760 473.700 88.020 ;
        RECT 821.660 87.760 821.920 88.020 ;
        RECT 821.660 19.080 821.920 19.340 ;
        RECT 827.640 19.080 827.900 19.340 ;
      LAYER met2 ;
        RECT 406.740 749.710 407.000 750.030 ;
        RECT 406.800 482.110 406.940 749.710 ;
        RECT 467.920 749.090 468.180 749.350 ;
        RECT 468.630 749.090 468.910 750.000 ;
        RECT 467.920 749.030 468.910 749.090 ;
        RECT 467.980 748.950 468.910 749.030 ;
        RECT 468.630 746.000 468.910 748.950 ;
        RECT 471.850 500.000 472.130 504.000 ;
        RECT 471.890 499.790 472.030 500.000 ;
        RECT 471.830 499.470 472.090 499.790 ;
        RECT 471.140 497.430 471.400 497.750 ;
        RECT 471.200 482.110 471.340 497.430 ;
        RECT 406.740 481.790 407.000 482.110 ;
        RECT 471.140 481.790 471.400 482.110 ;
        RECT 473.440 481.790 473.700 482.110 ;
        RECT 473.500 88.050 473.640 481.790 ;
        RECT 473.440 87.730 473.700 88.050 ;
        RECT 821.660 87.730 821.920 88.050 ;
        RECT 821.720 19.370 821.860 87.730 ;
        RECT 821.660 19.050 821.920 19.370 ;
        RECT 827.640 19.050 827.900 19.370 ;
        RECT 827.700 2.400 827.840 19.050 ;
        RECT 827.490 -4.800 828.050 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.960 499.700 585.280 499.760 ;
        RECT 584.960 499.500 585.420 499.700 ;
        RECT 585.280 497.320 585.420 499.500 ;
        RECT 586.110 497.320 586.430 497.380 ;
        RECT 585.280 497.180 586.430 497.320 ;
        RECT 586.110 497.120 586.430 497.180 ;
      LAYER via ;
        RECT 584.990 499.500 585.250 499.760 ;
        RECT 586.140 497.120 586.400 497.380 ;
      LAYER met2 ;
        RECT 585.010 500.000 585.290 504.000 ;
        RECT 585.050 499.790 585.190 500.000 ;
        RECT 584.990 499.470 585.250 499.790 ;
        RECT 586.130 497.235 586.410 497.605 ;
        RECT 586.140 497.090 586.400 497.235 ;
        RECT 2180.490 453.035 2180.770 453.405 ;
        RECT 2180.560 82.870 2180.700 453.035 ;
        RECT 2180.560 82.730 2185.760 82.870 ;
        RECT 2185.620 2.400 2185.760 82.730 ;
        RECT 2185.410 -4.800 2185.970 2.400 ;
      LAYER via2 ;
        RECT 586.130 497.280 586.410 497.560 ;
        RECT 2180.490 453.080 2180.770 453.360 ;
      LAYER met3 ;
        RECT 586.105 497.580 586.435 497.585 ;
        RECT 586.105 497.570 586.690 497.580 ;
        RECT 586.105 497.270 586.890 497.570 ;
        RECT 586.105 497.260 586.690 497.270 ;
        RECT 586.105 497.255 586.435 497.260 ;
        RECT 586.310 453.370 586.690 453.380 ;
        RECT 2180.465 453.370 2180.795 453.385 ;
        RECT 586.310 453.070 2180.795 453.370 ;
        RECT 586.310 453.060 586.690 453.070 ;
        RECT 2180.465 453.055 2180.795 453.070 ;
      LAYER via3 ;
        RECT 586.340 497.260 586.660 497.580 ;
        RECT 586.340 453.060 586.660 453.380 ;
      LAYER met4 ;
        RECT 586.335 497.255 586.665 497.585 ;
        RECT 586.350 453.385 586.650 497.255 ;
        RECT 586.335 453.055 586.665 453.385 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.340 499.160 586.660 499.420 ;
        RECT 586.430 497.660 586.570 499.160 ;
        RECT 587.490 497.660 587.810 497.720 ;
        RECT 586.430 497.520 587.810 497.660 ;
        RECT 587.490 497.460 587.810 497.520 ;
        RECT 587.490 480.660 587.810 480.720 ;
        RECT 588.410 480.660 588.730 480.720 ;
        RECT 587.490 480.520 588.730 480.660 ;
        RECT 587.490 480.460 587.810 480.520 ;
        RECT 588.410 480.460 588.730 480.520 ;
        RECT 588.410 424.220 588.730 424.280 ;
        RECT 2201.170 424.220 2201.490 424.280 ;
        RECT 588.410 424.080 2201.490 424.220 ;
        RECT 588.410 424.020 588.730 424.080 ;
        RECT 2201.170 424.020 2201.490 424.080 ;
      LAYER via ;
        RECT 586.370 499.160 586.630 499.420 ;
        RECT 587.520 497.460 587.780 497.720 ;
        RECT 587.520 480.460 587.780 480.720 ;
        RECT 588.440 480.460 588.700 480.720 ;
        RECT 588.440 424.020 588.700 424.280 ;
        RECT 2201.200 424.020 2201.460 424.280 ;
      LAYER met2 ;
        RECT 586.390 500.000 586.670 504.000 ;
        RECT 586.430 499.450 586.570 500.000 ;
        RECT 586.370 499.130 586.630 499.450 ;
        RECT 587.520 497.430 587.780 497.750 ;
        RECT 587.580 480.750 587.720 497.430 ;
        RECT 587.520 480.430 587.780 480.750 ;
        RECT 588.440 480.430 588.700 480.750 ;
        RECT 588.500 424.310 588.640 480.430 ;
        RECT 588.440 423.990 588.700 424.310 ;
        RECT 2201.200 423.990 2201.460 424.310 ;
        RECT 2201.260 17.410 2201.400 423.990 ;
        RECT 2201.260 17.270 2202.320 17.410 ;
        RECT 2202.180 2.400 2202.320 17.270 ;
        RECT 2201.970 -4.800 2202.530 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 585.740 500.240 587.950 500.380 ;
        RECT 585.740 498.400 585.880 500.240 ;
        RECT 587.810 499.760 587.950 500.240 ;
        RECT 587.720 499.500 588.040 499.760 ;
        RECT 585.650 498.140 585.970 498.400 ;
        RECT 585.650 491.540 585.970 491.600 ;
        RECT 587.950 491.540 588.270 491.600 ;
        RECT 585.650 491.400 588.270 491.540 ;
        RECT 585.650 491.340 585.970 491.400 ;
        RECT 587.950 491.340 588.270 491.400 ;
        RECT 587.950 197.780 588.270 197.840 ;
        RECT 2214.970 197.780 2215.290 197.840 ;
        RECT 587.950 197.640 2215.290 197.780 ;
        RECT 587.950 197.580 588.270 197.640 ;
        RECT 2214.970 197.580 2215.290 197.640 ;
      LAYER via ;
        RECT 587.750 499.500 588.010 499.760 ;
        RECT 585.680 498.140 585.940 498.400 ;
        RECT 585.680 491.340 585.940 491.600 ;
        RECT 587.980 491.340 588.240 491.600 ;
        RECT 587.980 197.580 588.240 197.840 ;
        RECT 2215.000 197.580 2215.260 197.840 ;
      LAYER met2 ;
        RECT 587.770 500.000 588.050 504.000 ;
        RECT 587.810 499.790 587.950 500.000 ;
        RECT 587.750 499.470 588.010 499.790 ;
        RECT 585.680 498.110 585.940 498.430 ;
        RECT 585.740 491.630 585.880 498.110 ;
        RECT 585.680 491.310 585.940 491.630 ;
        RECT 587.980 491.310 588.240 491.630 ;
        RECT 588.040 474.880 588.180 491.310 ;
        RECT 587.580 474.740 588.180 474.880 ;
        RECT 587.580 473.690 587.720 474.740 ;
        RECT 587.580 473.550 588.180 473.690 ;
        RECT 588.040 197.870 588.180 473.550 ;
        RECT 587.980 197.550 588.240 197.870 ;
        RECT 2215.000 197.550 2215.260 197.870 ;
        RECT 2215.060 82.870 2215.200 197.550 ;
        RECT 2215.060 82.730 2218.880 82.870 ;
        RECT 2218.740 2.400 2218.880 82.730 ;
        RECT 2218.530 -4.800 2219.090 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 589.100 499.700 589.420 499.760 ;
        RECT 588.960 499.500 589.420 499.700 ;
        RECT 588.960 497.720 589.100 499.500 ;
        RECT 588.870 497.460 589.190 497.720 ;
        RECT 588.870 431.360 589.190 431.420 ;
        RECT 2229.230 431.360 2229.550 431.420 ;
        RECT 588.870 431.220 2229.550 431.360 ;
        RECT 588.870 431.160 589.190 431.220 ;
        RECT 2229.230 431.160 2229.550 431.220 ;
        RECT 2229.230 18.940 2229.550 19.000 ;
        RECT 2235.210 18.940 2235.530 19.000 ;
        RECT 2229.230 18.800 2235.530 18.940 ;
        RECT 2229.230 18.740 2229.550 18.800 ;
        RECT 2235.210 18.740 2235.530 18.800 ;
      LAYER via ;
        RECT 589.130 499.500 589.390 499.760 ;
        RECT 588.900 497.460 589.160 497.720 ;
        RECT 588.900 431.160 589.160 431.420 ;
        RECT 2229.260 431.160 2229.520 431.420 ;
        RECT 2229.260 18.740 2229.520 19.000 ;
        RECT 2235.240 18.740 2235.500 19.000 ;
      LAYER met2 ;
        RECT 589.150 500.000 589.430 504.000 ;
        RECT 589.190 499.790 589.330 500.000 ;
        RECT 589.130 499.470 589.390 499.790 ;
        RECT 588.900 497.430 589.160 497.750 ;
        RECT 588.960 431.450 589.100 497.430 ;
        RECT 588.900 431.130 589.160 431.450 ;
        RECT 2229.260 431.130 2229.520 431.450 ;
        RECT 2229.320 19.030 2229.460 431.130 ;
        RECT 2229.260 18.710 2229.520 19.030 ;
        RECT 2235.240 18.710 2235.500 19.030 ;
        RECT 2235.300 2.400 2235.440 18.710 ;
        RECT 2235.090 -4.800 2235.650 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.530 500.000 590.810 504.000 ;
        RECT 590.570 498.680 590.710 500.000 ;
        RECT 590.570 498.540 590.940 498.680 ;
        RECT 590.800 498.000 590.940 498.540 ;
        RECT 590.800 497.860 591.400 498.000 ;
        RECT 591.260 485.365 591.400 497.860 ;
        RECT 591.190 484.995 591.470 485.365 ;
        RECT 2249.490 87.195 2249.770 87.565 ;
        RECT 2249.560 82.870 2249.700 87.195 ;
        RECT 2249.560 82.730 2252.000 82.870 ;
        RECT 2251.860 2.400 2252.000 82.730 ;
        RECT 2251.650 -4.800 2252.210 2.400 ;
      LAYER via2 ;
        RECT 591.190 485.040 591.470 485.320 ;
        RECT 2249.490 87.240 2249.770 87.520 ;
      LAYER met3 ;
        RECT 591.165 485.330 591.495 485.345 ;
        RECT 591.830 485.330 592.210 485.340 ;
        RECT 591.165 485.030 592.210 485.330 ;
        RECT 591.165 485.015 591.495 485.030 ;
        RECT 591.830 485.020 592.210 485.030 ;
        RECT 591.830 87.530 592.210 87.540 ;
        RECT 2249.465 87.530 2249.795 87.545 ;
        RECT 591.830 87.230 2249.795 87.530 ;
        RECT 591.830 87.220 592.210 87.230 ;
        RECT 2249.465 87.215 2249.795 87.230 ;
      LAYER via3 ;
        RECT 591.860 485.020 592.180 485.340 ;
        RECT 591.860 87.220 592.180 87.540 ;
      LAYER met4 ;
        RECT 591.855 485.015 592.185 485.345 ;
        RECT 591.870 87.545 592.170 485.015 ;
        RECT 591.855 87.215 592.185 87.545 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 591.860 499.500 592.180 499.760 ;
        RECT 591.950 498.060 592.090 499.500 ;
        RECT 591.950 497.860 592.410 498.060 ;
        RECT 592.090 497.800 592.410 497.860 ;
      LAYER via ;
        RECT 591.890 499.500 592.150 499.760 ;
        RECT 592.120 497.800 592.380 498.060 ;
      LAYER met2 ;
        RECT 591.910 500.000 592.190 504.000 ;
        RECT 591.950 499.790 592.090 500.000 ;
        RECT 591.890 499.470 592.150 499.790 ;
        RECT 592.120 497.770 592.380 498.090 ;
        RECT 592.180 486.045 592.320 497.770 ;
        RECT 592.110 485.675 592.390 486.045 ;
        RECT 2263.290 86.515 2263.570 86.885 ;
        RECT 2263.360 82.870 2263.500 86.515 ;
        RECT 2263.360 82.730 2268.560 82.870 ;
        RECT 2268.420 2.400 2268.560 82.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
      LAYER via2 ;
        RECT 592.110 485.720 592.390 486.000 ;
        RECT 2263.290 86.560 2263.570 86.840 ;
      LAYER met3 ;
        RECT 592.085 486.010 592.415 486.025 ;
        RECT 592.750 486.010 593.130 486.020 ;
        RECT 592.085 485.710 593.130 486.010 ;
        RECT 592.085 485.695 592.415 485.710 ;
        RECT 592.750 485.700 593.130 485.710 ;
        RECT 592.750 86.850 593.130 86.860 ;
        RECT 2263.265 86.850 2263.595 86.865 ;
        RECT 592.750 86.550 2263.595 86.850 ;
        RECT 592.750 86.540 593.130 86.550 ;
        RECT 2263.265 86.535 2263.595 86.550 ;
      LAYER via3 ;
        RECT 592.780 485.700 593.100 486.020 ;
        RECT 592.780 86.540 593.100 86.860 ;
      LAYER met4 ;
        RECT 592.775 485.695 593.105 486.025 ;
        RECT 592.790 86.865 593.090 485.695 ;
        RECT 592.775 86.535 593.105 86.865 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.240 499.700 593.560 499.760 ;
        RECT 593.240 499.560 595.080 499.700 ;
        RECT 593.240 499.500 593.560 499.560 ;
        RECT 594.940 498.060 595.080 499.560 ;
        RECT 594.850 497.800 595.170 498.060 ;
        RECT 594.850 487.120 595.170 487.180 ;
        RECT 596.690 487.120 597.010 487.180 ;
        RECT 594.850 486.980 597.010 487.120 ;
        RECT 594.850 486.920 595.170 486.980 ;
        RECT 596.690 486.920 597.010 486.980 ;
        RECT 596.690 459.240 597.010 459.300 ;
        RECT 2283.970 459.240 2284.290 459.300 ;
        RECT 596.690 459.100 2284.290 459.240 ;
        RECT 596.690 459.040 597.010 459.100 ;
        RECT 2283.970 459.040 2284.290 459.100 ;
      LAYER via ;
        RECT 593.270 499.500 593.530 499.760 ;
        RECT 594.880 497.800 595.140 498.060 ;
        RECT 594.880 486.920 595.140 487.180 ;
        RECT 596.720 486.920 596.980 487.180 ;
        RECT 596.720 459.040 596.980 459.300 ;
        RECT 2284.000 459.040 2284.260 459.300 ;
      LAYER met2 ;
        RECT 593.290 500.000 593.570 504.000 ;
        RECT 593.330 499.790 593.470 500.000 ;
        RECT 593.270 499.470 593.530 499.790 ;
        RECT 594.880 497.770 595.140 498.090 ;
        RECT 594.940 487.210 595.080 497.770 ;
        RECT 594.880 486.890 595.140 487.210 ;
        RECT 596.720 486.890 596.980 487.210 ;
        RECT 596.780 459.330 596.920 486.890 ;
        RECT 596.720 459.010 596.980 459.330 ;
        RECT 2284.000 459.010 2284.260 459.330 ;
        RECT 2284.060 17.410 2284.200 459.010 ;
        RECT 2284.060 17.270 2285.120 17.410 ;
        RECT 2284.980 2.400 2285.120 17.270 ;
        RECT 2284.770 -4.800 2285.330 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 87.620 593.790 87.680 ;
        RECT 2297.770 87.620 2298.090 87.680 ;
        RECT 593.470 87.480 2298.090 87.620 ;
        RECT 593.470 87.420 593.790 87.480 ;
        RECT 2297.770 87.420 2298.090 87.480 ;
      LAYER via ;
        RECT 593.500 87.420 593.760 87.680 ;
        RECT 2297.800 87.420 2298.060 87.680 ;
      LAYER met2 ;
        RECT 594.670 500.000 594.950 504.000 ;
        RECT 594.710 499.815 594.850 500.000 ;
        RECT 594.640 499.445 594.920 499.815 ;
        RECT 593.490 497.915 593.770 498.285 ;
        RECT 593.560 87.710 593.700 497.915 ;
        RECT 593.500 87.390 593.760 87.710 ;
        RECT 2297.800 87.390 2298.060 87.710 ;
        RECT 2297.860 82.870 2298.000 87.390 ;
        RECT 2297.860 82.730 2301.680 82.870 ;
        RECT 2301.540 2.400 2301.680 82.730 ;
        RECT 2301.330 -4.800 2301.890 2.400 ;
      LAYER via2 ;
        RECT 594.640 499.490 594.920 499.770 ;
        RECT 593.490 497.960 593.770 498.240 ;
      LAYER met3 ;
        RECT 594.615 499.465 594.945 499.795 ;
        RECT 594.630 498.930 594.930 499.465 ;
        RECT 593.710 498.630 594.930 498.930 ;
        RECT 593.710 498.265 594.010 498.630 ;
        RECT 593.465 497.950 594.010 498.265 ;
        RECT 593.465 497.935 593.795 497.950 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.000 499.500 596.320 499.760 ;
        RECT 596.090 498.000 596.230 499.500 ;
        RECT 596.090 497.860 597.380 498.000 ;
        RECT 597.240 497.380 597.380 497.860 ;
        RECT 597.150 497.120 597.470 497.380 ;
        RECT 593.930 484.060 594.250 484.120 ;
        RECT 597.150 484.060 597.470 484.120 ;
        RECT 593.930 483.920 597.470 484.060 ;
        RECT 593.930 483.860 594.250 483.920 ;
        RECT 597.150 483.860 597.470 483.920 ;
        RECT 593.930 87.280 594.250 87.340 ;
        RECT 2312.030 87.280 2312.350 87.340 ;
        RECT 593.930 87.140 2312.350 87.280 ;
        RECT 593.930 87.080 594.250 87.140 ;
        RECT 2312.030 87.080 2312.350 87.140 ;
        RECT 2312.030 18.600 2312.350 18.660 ;
        RECT 2318.010 18.600 2318.330 18.660 ;
        RECT 2312.030 18.460 2318.330 18.600 ;
        RECT 2312.030 18.400 2312.350 18.460 ;
        RECT 2318.010 18.400 2318.330 18.460 ;
      LAYER via ;
        RECT 596.030 499.500 596.290 499.760 ;
        RECT 597.180 497.120 597.440 497.380 ;
        RECT 593.960 483.860 594.220 484.120 ;
        RECT 597.180 483.860 597.440 484.120 ;
        RECT 593.960 87.080 594.220 87.340 ;
        RECT 2312.060 87.080 2312.320 87.340 ;
        RECT 2312.060 18.400 2312.320 18.660 ;
        RECT 2318.040 18.400 2318.300 18.660 ;
      LAYER met2 ;
        RECT 596.050 500.000 596.330 504.000 ;
        RECT 596.090 499.790 596.230 500.000 ;
        RECT 596.030 499.470 596.290 499.790 ;
        RECT 597.180 497.090 597.440 497.410 ;
        RECT 597.240 484.150 597.380 497.090 ;
        RECT 593.960 483.830 594.220 484.150 ;
        RECT 597.180 483.830 597.440 484.150 ;
        RECT 594.020 87.370 594.160 483.830 ;
        RECT 593.960 87.050 594.220 87.370 ;
        RECT 2312.060 87.050 2312.320 87.370 ;
        RECT 2312.120 18.690 2312.260 87.050 ;
        RECT 2312.060 18.370 2312.320 18.690 ;
        RECT 2318.040 18.370 2318.300 18.690 ;
        RECT 2318.100 2.400 2318.240 18.370 ;
        RECT 2317.890 -4.800 2318.450 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 597.380 499.500 597.700 499.760 ;
        RECT 597.470 499.080 597.610 499.500 ;
        RECT 597.470 498.880 597.930 499.080 ;
        RECT 597.610 498.820 597.930 498.880 ;
        RECT 594.390 483.040 594.710 483.100 ;
        RECT 598.070 483.040 598.390 483.100 ;
        RECT 594.390 482.900 598.390 483.040 ;
        RECT 594.390 482.840 594.710 482.900 ;
        RECT 598.070 482.840 598.390 482.900 ;
        RECT 594.390 94.080 594.710 94.140 ;
        RECT 2332.270 94.080 2332.590 94.140 ;
        RECT 594.390 93.940 2332.590 94.080 ;
        RECT 594.390 93.880 594.710 93.940 ;
        RECT 2332.270 93.880 2332.590 93.940 ;
      LAYER via ;
        RECT 597.410 499.500 597.670 499.760 ;
        RECT 597.640 498.820 597.900 499.080 ;
        RECT 594.420 482.840 594.680 483.100 ;
        RECT 598.100 482.840 598.360 483.100 ;
        RECT 594.420 93.880 594.680 94.140 ;
        RECT 2332.300 93.880 2332.560 94.140 ;
      LAYER met2 ;
        RECT 597.430 500.000 597.710 504.000 ;
        RECT 597.470 499.790 597.610 500.000 ;
        RECT 597.410 499.470 597.670 499.790 ;
        RECT 597.640 498.790 597.900 499.110 ;
        RECT 597.700 485.080 597.840 498.790 ;
        RECT 597.700 484.940 598.300 485.080 ;
        RECT 598.160 483.130 598.300 484.940 ;
        RECT 594.420 482.810 594.680 483.130 ;
        RECT 598.100 482.810 598.360 483.130 ;
        RECT 594.480 94.170 594.620 482.810 ;
        RECT 594.420 93.850 594.680 94.170 ;
        RECT 2332.300 93.850 2332.560 94.170 ;
        RECT 2332.360 82.870 2332.500 93.850 ;
        RECT 2332.360 82.730 2334.800 82.870 ;
        RECT 2334.660 2.400 2334.800 82.730 ;
        RECT 2334.450 -4.800 2335.010 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 404.410 762.520 404.730 762.580 ;
        RECT 473.410 762.520 473.730 762.580 ;
        RECT 404.410 762.380 473.730 762.520 ;
        RECT 404.410 762.320 404.730 762.380 ;
        RECT 473.410 762.320 473.730 762.380 ;
        RECT 404.410 501.060 404.730 501.120 ;
        RECT 404.410 500.920 434.770 501.060 ;
        RECT 404.410 500.860 404.730 500.920 ;
        RECT 434.630 500.720 434.770 500.920 ;
        RECT 434.630 500.580 469.270 500.720 ;
        RECT 469.130 500.380 469.270 500.580 ;
        RECT 469.130 500.240 473.410 500.380 ;
        RECT 470.510 497.720 470.650 500.240 ;
        RECT 473.270 499.760 473.410 500.240 ;
        RECT 473.180 499.500 473.500 499.760 ;
        RECT 470.190 497.520 470.650 497.720 ;
        RECT 470.190 497.460 470.510 497.520 ;
        RECT 469.270 472.840 469.590 472.900 ;
        RECT 470.190 472.840 470.510 472.900 ;
        RECT 469.270 472.700 470.510 472.840 ;
        RECT 469.270 472.640 469.590 472.700 ;
        RECT 470.190 472.640 470.510 472.700 ;
        RECT 469.270 94.760 469.590 94.820 ;
        RECT 841.870 94.760 842.190 94.820 ;
        RECT 469.270 94.620 842.190 94.760 ;
        RECT 469.270 94.560 469.590 94.620 ;
        RECT 841.870 94.560 842.190 94.620 ;
      LAYER via ;
        RECT 404.440 762.320 404.700 762.580 ;
        RECT 473.440 762.320 473.700 762.580 ;
        RECT 404.440 500.860 404.700 501.120 ;
        RECT 473.210 499.500 473.470 499.760 ;
        RECT 470.220 497.460 470.480 497.720 ;
        RECT 469.300 472.640 469.560 472.900 ;
        RECT 470.220 472.640 470.480 472.900 ;
        RECT 469.300 94.560 469.560 94.820 ;
        RECT 841.900 94.560 842.160 94.820 ;
      LAYER met2 ;
        RECT 404.440 762.290 404.700 762.610 ;
        RECT 473.440 762.290 473.700 762.610 ;
        RECT 404.500 501.150 404.640 762.290 ;
        RECT 473.500 749.770 473.640 762.290 ;
        RECT 474.150 749.770 474.430 750.000 ;
        RECT 473.500 749.630 474.430 749.770 ;
        RECT 474.150 746.000 474.430 749.630 ;
        RECT 404.440 500.830 404.700 501.150 ;
        RECT 473.230 500.000 473.510 504.000 ;
        RECT 473.270 499.790 473.410 500.000 ;
        RECT 473.210 499.470 473.470 499.790 ;
        RECT 470.220 497.430 470.480 497.750 ;
        RECT 470.280 472.930 470.420 497.430 ;
        RECT 469.300 472.610 469.560 472.930 ;
        RECT 470.220 472.610 470.480 472.930 ;
        RECT 469.360 94.850 469.500 472.610 ;
        RECT 469.300 94.530 469.560 94.850 ;
        RECT 841.900 94.530 842.160 94.850 ;
        RECT 841.960 82.870 842.100 94.530 ;
        RECT 841.960 82.730 844.400 82.870 ;
        RECT 844.260 2.400 844.400 82.730 ;
        RECT 844.050 -4.800 844.610 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.270 500.000 461.550 504.000 ;
        RECT 461.310 499.815 461.450 500.000 ;
        RECT 461.240 499.445 461.520 499.815 ;
        RECT 696.990 94.675 697.270 95.045 ;
        RECT 697.060 82.870 697.200 94.675 ;
        RECT 697.060 82.730 700.880 82.870 ;
        RECT 700.740 2.400 700.880 82.730 ;
        RECT 700.530 -4.800 701.090 2.400 ;
      LAYER via2 ;
        RECT 461.240 499.490 461.520 499.770 ;
        RECT 696.990 94.720 697.270 95.000 ;
      LAYER met3 ;
        RECT 461.215 499.465 461.545 499.795 ;
        RECT 457.510 498.250 457.890 498.260 ;
        RECT 461.230 498.250 461.530 499.465 ;
        RECT 457.510 497.950 461.530 498.250 ;
        RECT 457.510 497.940 457.890 497.950 ;
        RECT 457.510 95.010 457.890 95.020 ;
        RECT 696.965 95.010 697.295 95.025 ;
        RECT 457.510 94.710 697.295 95.010 ;
        RECT 457.510 94.700 457.890 94.710 ;
        RECT 696.965 94.695 697.295 94.710 ;
      LAYER via3 ;
        RECT 457.540 497.940 457.860 498.260 ;
        RECT 457.540 94.700 457.860 95.020 ;
      LAYER met4 ;
        RECT 457.535 497.935 457.865 498.265 ;
        RECT 457.550 95.025 457.850 497.935 ;
        RECT 457.535 94.695 457.865 95.025 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 599.220 499.360 599.540 499.420 ;
        RECT 599.080 499.160 599.540 499.360 ;
        RECT 599.080 498.740 599.220 499.160 ;
        RECT 598.990 498.480 599.310 498.740 ;
      LAYER via ;
        RECT 599.250 499.160 599.510 499.420 ;
        RECT 599.020 498.480 599.280 498.740 ;
      LAYER met2 ;
        RECT 599.270 500.000 599.550 504.000 ;
        RECT 599.310 499.450 599.450 500.000 ;
        RECT 599.250 499.130 599.510 499.450 ;
        RECT 599.020 498.450 599.280 498.770 ;
        RECT 599.080 486.045 599.220 498.450 ;
        RECT 599.010 485.675 599.290 486.045 ;
        RECT 2352.990 93.995 2353.270 94.365 ;
        RECT 2353.060 82.870 2353.200 93.995 ;
        RECT 2353.060 82.730 2356.880 82.870 ;
        RECT 2356.740 2.400 2356.880 82.730 ;
        RECT 2356.530 -4.800 2357.090 2.400 ;
      LAYER via2 ;
        RECT 599.010 485.720 599.290 486.000 ;
        RECT 2352.990 94.040 2353.270 94.320 ;
      LAYER met3 ;
        RECT 598.985 486.020 599.315 486.025 ;
        RECT 598.985 486.010 599.570 486.020 ;
        RECT 598.985 485.710 599.770 486.010 ;
        RECT 598.985 485.700 599.570 485.710 ;
        RECT 598.985 485.695 599.315 485.700 ;
        RECT 599.190 94.330 599.570 94.340 ;
        RECT 2352.965 94.330 2353.295 94.345 ;
        RECT 599.190 94.030 2353.295 94.330 ;
        RECT 599.190 94.020 599.570 94.030 ;
        RECT 2352.965 94.015 2353.295 94.030 ;
      LAYER via3 ;
        RECT 599.220 485.700 599.540 486.020 ;
        RECT 599.220 94.020 599.540 94.340 ;
      LAYER met4 ;
        RECT 599.215 485.695 599.545 486.025 ;
        RECT 599.230 94.345 599.530 485.695 ;
        RECT 599.215 94.015 599.545 94.345 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.600 499.500 600.920 499.760 ;
        RECT 600.690 498.340 600.830 499.500 ;
        RECT 604.050 498.340 604.370 498.400 ;
        RECT 600.690 498.200 604.370 498.340 ;
        RECT 604.050 498.140 604.370 498.200 ;
        RECT 604.510 451.760 604.830 451.820 ;
        RECT 2367.230 451.760 2367.550 451.820 ;
        RECT 604.510 451.620 2367.550 451.760 ;
        RECT 604.510 451.560 604.830 451.620 ;
        RECT 2367.230 451.560 2367.550 451.620 ;
        RECT 2367.230 17.920 2367.550 17.980 ;
        RECT 2373.210 17.920 2373.530 17.980 ;
        RECT 2367.230 17.780 2373.530 17.920 ;
        RECT 2367.230 17.720 2367.550 17.780 ;
        RECT 2373.210 17.720 2373.530 17.780 ;
      LAYER via ;
        RECT 600.630 499.500 600.890 499.760 ;
        RECT 604.080 498.140 604.340 498.400 ;
        RECT 604.540 451.560 604.800 451.820 ;
        RECT 2367.260 451.560 2367.520 451.820 ;
        RECT 2367.260 17.720 2367.520 17.980 ;
        RECT 2373.240 17.720 2373.500 17.980 ;
      LAYER met2 ;
        RECT 600.650 500.000 600.930 504.000 ;
        RECT 600.690 499.790 600.830 500.000 ;
        RECT 600.630 499.470 600.890 499.790 ;
        RECT 604.080 498.110 604.340 498.430 ;
        RECT 604.140 485.250 604.280 498.110 ;
        RECT 604.140 485.110 604.740 485.250 ;
        RECT 604.600 451.850 604.740 485.110 ;
        RECT 604.540 451.530 604.800 451.850 ;
        RECT 2367.260 451.530 2367.520 451.850 ;
        RECT 2367.320 18.010 2367.460 451.530 ;
        RECT 2367.260 17.690 2367.520 18.010 ;
        RECT 2373.240 17.690 2373.500 18.010 ;
        RECT 2373.300 2.400 2373.440 17.690 ;
        RECT 2373.090 -4.800 2373.650 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 602.210 93.740 602.530 93.800 ;
        RECT 2387.470 93.740 2387.790 93.800 ;
        RECT 602.210 93.600 2387.790 93.740 ;
        RECT 602.210 93.540 602.530 93.600 ;
        RECT 2387.470 93.540 2387.790 93.600 ;
      LAYER via ;
        RECT 602.240 93.540 602.500 93.800 ;
        RECT 2387.500 93.540 2387.760 93.800 ;
      LAYER met2 ;
        RECT 602.030 500.000 602.310 504.000 ;
        RECT 602.070 499.815 602.210 500.000 ;
        RECT 602.000 499.445 602.280 499.815 ;
        RECT 602.230 497.235 602.510 497.605 ;
        RECT 602.300 93.830 602.440 497.235 ;
        RECT 602.240 93.510 602.500 93.830 ;
        RECT 2387.500 93.510 2387.760 93.830 ;
        RECT 2387.560 82.870 2387.700 93.510 ;
        RECT 2387.560 82.730 2390.000 82.870 ;
        RECT 2389.860 2.400 2390.000 82.730 ;
        RECT 2389.650 -4.800 2390.210 2.400 ;
      LAYER via2 ;
        RECT 602.000 499.490 602.280 499.770 ;
        RECT 602.230 497.280 602.510 497.560 ;
      LAYER met3 ;
        RECT 601.975 499.465 602.305 499.795 ;
        RECT 601.990 497.585 602.290 499.465 ;
        RECT 601.990 497.270 602.535 497.585 ;
        RECT 602.205 497.255 602.535 497.270 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 603.360 499.500 603.680 499.760 ;
        RECT 603.450 499.360 603.590 499.500 ;
        RECT 603.450 499.220 603.820 499.360 ;
        RECT 603.680 499.080 603.820 499.220 ;
        RECT 603.590 498.820 603.910 499.080 ;
        RECT 600.370 486.780 600.690 486.840 ;
        RECT 603.590 486.780 603.910 486.840 ;
        RECT 600.370 486.640 603.910 486.780 ;
        RECT 600.370 486.580 600.690 486.640 ;
        RECT 603.590 486.580 603.910 486.640 ;
        RECT 600.830 25.740 601.150 25.800 ;
        RECT 2406.330 25.740 2406.650 25.800 ;
        RECT 600.830 25.600 2406.650 25.740 ;
        RECT 600.830 25.540 601.150 25.600 ;
        RECT 2406.330 25.540 2406.650 25.600 ;
      LAYER via ;
        RECT 603.390 499.500 603.650 499.760 ;
        RECT 603.620 498.820 603.880 499.080 ;
        RECT 600.400 486.580 600.660 486.840 ;
        RECT 603.620 486.580 603.880 486.840 ;
        RECT 600.860 25.540 601.120 25.800 ;
        RECT 2406.360 25.540 2406.620 25.800 ;
      LAYER met2 ;
        RECT 603.410 500.000 603.690 504.000 ;
        RECT 603.450 499.790 603.590 500.000 ;
        RECT 603.390 499.470 603.650 499.790 ;
        RECT 603.620 498.790 603.880 499.110 ;
        RECT 603.680 486.870 603.820 498.790 ;
        RECT 600.400 486.550 600.660 486.870 ;
        RECT 603.620 486.550 603.880 486.870 ;
        RECT 600.460 448.570 600.600 486.550 ;
        RECT 600.460 448.430 601.060 448.570 ;
        RECT 600.920 25.830 601.060 448.430 ;
        RECT 600.860 25.510 601.120 25.830 ;
        RECT 2406.360 25.510 2406.620 25.830 ;
        RECT 2406.420 2.400 2406.560 25.510 ;
        RECT 2406.210 -4.800 2406.770 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 604.740 499.500 605.060 499.760 ;
        RECT 604.830 497.380 604.970 499.500 ;
        RECT 604.830 497.180 605.290 497.380 ;
        RECT 604.970 497.120 605.290 497.180 ;
      LAYER via ;
        RECT 604.770 499.500 605.030 499.760 ;
        RECT 605.000 497.120 605.260 497.380 ;
      LAYER met2 ;
        RECT 604.790 500.000 605.070 504.000 ;
        RECT 604.830 499.790 604.970 500.000 ;
        RECT 604.770 499.470 605.030 499.790 ;
        RECT 605.000 497.090 605.260 497.410 ;
        RECT 605.060 486.725 605.200 497.090 ;
        RECT 604.990 486.355 605.270 486.725 ;
        RECT 2422.910 32.115 2423.190 32.485 ;
        RECT 2422.980 2.400 2423.120 32.115 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
      LAYER via2 ;
        RECT 604.990 486.400 605.270 486.680 ;
        RECT 2422.910 32.160 2423.190 32.440 ;
      LAYER met3 ;
        RECT 604.965 486.690 605.295 486.705 ;
        RECT 605.630 486.690 606.010 486.700 ;
        RECT 604.965 486.390 606.010 486.690 ;
        RECT 604.965 486.375 605.295 486.390 ;
        RECT 605.630 486.380 606.010 486.390 ;
        RECT 605.630 32.450 606.010 32.460 ;
        RECT 2422.885 32.450 2423.215 32.465 ;
        RECT 605.630 32.150 2423.215 32.450 ;
        RECT 605.630 32.140 606.010 32.150 ;
        RECT 2422.885 32.135 2423.215 32.150 ;
      LAYER via3 ;
        RECT 605.660 486.380 605.980 486.700 ;
        RECT 605.660 32.140 605.980 32.460 ;
      LAYER met4 ;
        RECT 605.655 486.375 605.985 486.705 ;
        RECT 605.670 32.465 605.970 486.375 ;
        RECT 605.655 32.135 605.985 32.465 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.120 498.820 606.440 499.080 ;
        RECT 606.210 498.400 606.350 498.820 ;
        RECT 605.890 498.200 606.350 498.400 ;
        RECT 605.890 498.140 606.210 498.200 ;
      LAYER via ;
        RECT 606.150 498.820 606.410 499.080 ;
        RECT 605.920 498.140 606.180 498.400 ;
      LAYER met2 ;
        RECT 606.170 500.000 606.450 504.000 ;
        RECT 606.210 499.110 606.350 500.000 ;
        RECT 606.150 498.790 606.410 499.110 ;
        RECT 605.920 498.110 606.180 498.430 ;
        RECT 605.980 484.685 606.120 498.110 ;
        RECT 605.910 484.315 606.190 484.685 ;
        RECT 2439.470 31.435 2439.750 31.805 ;
        RECT 2439.540 2.400 2439.680 31.435 ;
        RECT 2439.330 -4.800 2439.890 2.400 ;
      LAYER via2 ;
        RECT 605.910 484.360 606.190 484.640 ;
        RECT 2439.470 31.480 2439.750 31.760 ;
      LAYER met3 ;
        RECT 603.790 484.650 604.170 484.660 ;
        RECT 605.885 484.650 606.215 484.665 ;
        RECT 603.790 484.350 606.215 484.650 ;
        RECT 603.790 484.340 604.170 484.350 ;
        RECT 605.885 484.335 606.215 484.350 ;
        RECT 603.790 31.770 604.170 31.780 ;
        RECT 2439.445 31.770 2439.775 31.785 ;
        RECT 603.790 31.470 2439.775 31.770 ;
        RECT 603.790 31.460 604.170 31.470 ;
        RECT 2439.445 31.455 2439.775 31.470 ;
      LAYER via3 ;
        RECT 603.820 484.340 604.140 484.660 ;
        RECT 603.820 31.460 604.140 31.780 ;
      LAYER met4 ;
        RECT 603.815 484.335 604.145 484.665 ;
        RECT 603.830 31.785 604.130 484.335 ;
        RECT 603.815 31.455 604.145 31.785 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.490 101.900 610.810 101.960 ;
        RECT 2450.030 101.900 2450.350 101.960 ;
        RECT 610.490 101.760 2450.350 101.900 ;
        RECT 610.490 101.700 610.810 101.760 ;
        RECT 2450.030 101.700 2450.350 101.760 ;
        RECT 2450.030 17.580 2450.350 17.640 ;
        RECT 2456.010 17.580 2456.330 17.640 ;
        RECT 2450.030 17.440 2456.330 17.580 ;
        RECT 2450.030 17.380 2450.350 17.440 ;
        RECT 2456.010 17.380 2456.330 17.440 ;
      LAYER via ;
        RECT 610.520 101.700 610.780 101.960 ;
        RECT 2450.060 101.700 2450.320 101.960 ;
        RECT 2450.060 17.380 2450.320 17.640 ;
        RECT 2456.040 17.380 2456.300 17.640 ;
      LAYER met2 ;
        RECT 607.550 500.000 607.830 504.000 ;
        RECT 607.590 499.815 607.730 500.000 ;
        RECT 607.520 499.445 607.800 499.815 ;
        RECT 610.510 497.235 610.790 497.605 ;
        RECT 610.580 101.990 610.720 497.235 ;
        RECT 610.520 101.670 610.780 101.990 ;
        RECT 2450.060 101.670 2450.320 101.990 ;
        RECT 2450.120 17.670 2450.260 101.670 ;
        RECT 2450.060 17.350 2450.320 17.670 ;
        RECT 2456.040 17.350 2456.300 17.670 ;
        RECT 2456.100 2.400 2456.240 17.350 ;
        RECT 2455.890 -4.800 2456.450 2.400 ;
      LAYER via2 ;
        RECT 607.520 499.490 607.800 499.770 ;
        RECT 610.510 497.280 610.790 497.560 ;
      LAYER met3 ;
        RECT 607.495 499.465 607.825 499.795 ;
        RECT 607.510 497.570 607.810 499.465 ;
        RECT 610.485 497.570 610.815 497.585 ;
        RECT 607.510 497.270 610.815 497.570 ;
        RECT 610.485 497.255 610.815 497.270 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.030 101.560 610.350 101.620 ;
        RECT 2470.270 101.560 2470.590 101.620 ;
        RECT 610.030 101.420 2470.590 101.560 ;
        RECT 610.030 101.360 610.350 101.420 ;
        RECT 2470.270 101.360 2470.590 101.420 ;
      LAYER via ;
        RECT 610.060 101.360 610.320 101.620 ;
        RECT 2470.300 101.360 2470.560 101.620 ;
      LAYER met2 ;
        RECT 608.930 500.000 609.210 504.000 ;
        RECT 608.970 498.680 609.110 500.000 ;
        RECT 608.970 498.540 609.340 498.680 ;
        RECT 609.200 476.410 609.340 498.540 ;
        RECT 609.200 476.270 610.260 476.410 ;
        RECT 610.120 101.650 610.260 476.270 ;
        RECT 610.060 101.330 610.320 101.650 ;
        RECT 2470.300 101.330 2470.560 101.650 ;
        RECT 2470.360 82.870 2470.500 101.330 ;
        RECT 2470.360 82.730 2472.800 82.870 ;
        RECT 2472.660 2.400 2472.800 82.730 ;
        RECT 2472.450 -4.800 2473.010 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.950 101.220 611.270 101.280 ;
        RECT 2484.070 101.220 2484.390 101.280 ;
        RECT 610.950 101.080 2484.390 101.220 ;
        RECT 610.950 101.020 611.270 101.080 ;
        RECT 2484.070 101.020 2484.390 101.080 ;
      LAYER via ;
        RECT 610.980 101.020 611.240 101.280 ;
        RECT 2484.100 101.020 2484.360 101.280 ;
      LAYER met2 ;
        RECT 610.310 500.000 610.590 504.000 ;
        RECT 610.350 499.645 610.490 500.000 ;
        RECT 610.280 499.275 610.560 499.645 ;
        RECT 610.970 497.915 611.250 498.285 ;
        RECT 611.040 101.310 611.180 497.915 ;
        RECT 610.980 100.990 611.240 101.310 ;
        RECT 2484.100 100.990 2484.360 101.310 ;
        RECT 2484.160 82.870 2484.300 100.990 ;
        RECT 2484.160 82.730 2489.360 82.870 ;
        RECT 2489.220 2.400 2489.360 82.730 ;
        RECT 2489.010 -4.800 2489.570 2.400 ;
      LAYER via2 ;
        RECT 610.280 499.320 610.560 499.600 ;
        RECT 610.970 497.960 611.250 498.240 ;
      LAYER met3 ;
        RECT 610.255 499.610 610.585 499.625 ;
        RECT 610.255 499.310 611.260 499.610 ;
        RECT 610.255 499.295 610.585 499.310 ;
        RECT 610.960 498.265 611.260 499.310 ;
        RECT 610.945 497.935 611.275 498.265 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.640 499.700 611.960 499.760 ;
        RECT 611.640 499.560 613.250 499.700 ;
        RECT 611.640 499.500 611.960 499.560 ;
        RECT 611.410 498.000 611.730 498.060 ;
        RECT 613.110 498.000 613.250 499.560 ;
        RECT 611.410 497.860 613.250 498.000 ;
        RECT 611.410 497.800 611.730 497.860 ;
        RECT 609.570 472.160 609.890 472.220 ;
        RECT 611.410 472.160 611.730 472.220 ;
        RECT 609.570 472.020 611.730 472.160 ;
        RECT 609.570 471.960 609.890 472.020 ;
        RECT 611.410 471.960 611.730 472.020 ;
        RECT 609.570 100.880 609.890 100.940 ;
        RECT 2504.770 100.880 2505.090 100.940 ;
        RECT 609.570 100.740 2505.090 100.880 ;
        RECT 609.570 100.680 609.890 100.740 ;
        RECT 2504.770 100.680 2505.090 100.740 ;
      LAYER via ;
        RECT 611.670 499.500 611.930 499.760 ;
        RECT 611.440 497.800 611.700 498.060 ;
        RECT 609.600 471.960 609.860 472.220 ;
        RECT 611.440 471.960 611.700 472.220 ;
        RECT 609.600 100.680 609.860 100.940 ;
        RECT 2504.800 100.680 2505.060 100.940 ;
      LAYER met2 ;
        RECT 611.690 500.000 611.970 504.000 ;
        RECT 611.730 499.790 611.870 500.000 ;
        RECT 611.670 499.470 611.930 499.790 ;
        RECT 611.440 497.770 611.700 498.090 ;
        RECT 611.500 472.250 611.640 497.770 ;
        RECT 609.600 471.930 609.860 472.250 ;
        RECT 611.440 471.930 611.700 472.250 ;
        RECT 609.660 100.970 609.800 471.930 ;
        RECT 609.600 100.650 609.860 100.970 ;
        RECT 2504.800 100.650 2505.060 100.970 ;
        RECT 2504.860 17.410 2505.000 100.650 ;
        RECT 2504.860 17.270 2505.920 17.410 ;
        RECT 2505.780 2.400 2505.920 17.270 ;
        RECT 2505.570 -4.800 2506.130 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.070 500.000 475.350 504.000 ;
        RECT 475.110 498.965 475.250 500.000 ;
        RECT 475.040 498.595 475.320 498.965 ;
        RECT 862.590 100.115 862.870 100.485 ;
        RECT 862.660 82.870 862.800 100.115 ;
        RECT 862.660 82.730 866.480 82.870 ;
        RECT 866.340 2.400 866.480 82.730 ;
        RECT 866.130 -4.800 866.690 2.400 ;
      LAYER via2 ;
        RECT 475.040 498.640 475.320 498.920 ;
        RECT 862.590 100.160 862.870 100.440 ;
      LAYER met3 ;
        RECT 475.015 498.940 475.345 498.945 ;
        RECT 474.990 498.930 475.370 498.940 ;
        RECT 474.560 498.630 475.370 498.930 ;
        RECT 474.990 498.620 475.370 498.630 ;
        RECT 475.015 498.615 475.345 498.620 ;
        RECT 474.990 100.450 475.370 100.460 ;
        RECT 862.565 100.450 862.895 100.465 ;
        RECT 474.990 100.150 862.895 100.450 ;
        RECT 474.990 100.140 475.370 100.150 ;
        RECT 862.565 100.135 862.895 100.150 ;
      LAYER via3 ;
        RECT 475.020 498.620 475.340 498.940 ;
        RECT 475.020 100.140 475.340 100.460 ;
      LAYER met4 ;
        RECT 475.015 498.615 475.345 498.945 ;
        RECT 475.030 100.465 475.330 498.615 ;
        RECT 475.015 100.135 475.345 100.465 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.070 500.000 613.350 504.000 ;
        RECT 613.110 498.850 613.250 500.000 ;
        RECT 612.880 498.710 613.250 498.850 ;
        RECT 612.880 492.165 613.020 498.710 ;
        RECT 612.810 491.795 613.090 492.165 ;
        RECT 2522.270 30.755 2522.550 31.125 ;
        RECT 2522.340 2.400 2522.480 30.755 ;
        RECT 2522.130 -4.800 2522.690 2.400 ;
      LAYER via2 ;
        RECT 612.810 491.840 613.090 492.120 ;
        RECT 2522.270 30.800 2522.550 31.080 ;
      LAYER met3 ;
        RECT 610.230 492.130 610.610 492.140 ;
        RECT 612.785 492.130 613.115 492.145 ;
        RECT 610.230 491.830 613.115 492.130 ;
        RECT 610.230 491.820 610.610 491.830 ;
        RECT 612.785 491.815 613.115 491.830 ;
        RECT 610.230 31.090 610.610 31.100 ;
        RECT 2522.245 31.090 2522.575 31.105 ;
        RECT 610.230 30.790 2522.575 31.090 ;
        RECT 610.230 30.780 610.610 30.790 ;
        RECT 2522.245 30.775 2522.575 30.790 ;
      LAYER via3 ;
        RECT 610.260 491.820 610.580 492.140 ;
        RECT 610.260 30.780 610.580 31.100 ;
      LAYER met4 ;
        RECT 610.255 491.815 610.585 492.145 ;
        RECT 610.270 31.105 610.570 491.815 ;
        RECT 610.255 30.775 610.585 31.105 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.710 471.480 614.030 471.540 ;
        RECT 616.470 471.480 616.790 471.540 ;
        RECT 613.710 471.340 616.790 471.480 ;
        RECT 613.710 471.280 614.030 471.340 ;
        RECT 616.470 471.280 616.790 471.340 ;
        RECT 616.470 108.360 616.790 108.420 ;
        RECT 2532.830 108.360 2533.150 108.420 ;
        RECT 616.470 108.220 2533.150 108.360 ;
        RECT 616.470 108.160 616.790 108.220 ;
        RECT 2532.830 108.160 2533.150 108.220 ;
        RECT 2532.830 17.920 2533.150 17.980 ;
        RECT 2538.810 17.920 2539.130 17.980 ;
        RECT 2532.830 17.780 2539.130 17.920 ;
        RECT 2532.830 17.720 2533.150 17.780 ;
        RECT 2538.810 17.720 2539.130 17.780 ;
      LAYER via ;
        RECT 613.740 471.280 614.000 471.540 ;
        RECT 616.500 471.280 616.760 471.540 ;
        RECT 616.500 108.160 616.760 108.420 ;
        RECT 2532.860 108.160 2533.120 108.420 ;
        RECT 2532.860 17.720 2533.120 17.980 ;
        RECT 2538.840 17.720 2539.100 17.980 ;
      LAYER met2 ;
        RECT 614.450 500.000 614.730 504.000 ;
        RECT 614.490 498.850 614.630 500.000 ;
        RECT 614.260 498.710 614.630 498.850 ;
        RECT 614.260 473.690 614.400 498.710 ;
        RECT 613.800 473.550 614.400 473.690 ;
        RECT 613.800 471.570 613.940 473.550 ;
        RECT 613.740 471.250 614.000 471.570 ;
        RECT 616.500 471.250 616.760 471.570 ;
        RECT 616.560 108.450 616.700 471.250 ;
        RECT 616.500 108.130 616.760 108.450 ;
        RECT 2532.860 108.130 2533.120 108.450 ;
        RECT 2532.920 18.010 2533.060 108.130 ;
        RECT 2532.860 17.690 2533.120 18.010 ;
        RECT 2538.840 17.690 2539.100 18.010 ;
        RECT 2538.900 2.400 2539.040 17.690 ;
        RECT 2538.690 -4.800 2539.250 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.010 108.020 616.330 108.080 ;
        RECT 2553.070 108.020 2553.390 108.080 ;
        RECT 616.010 107.880 2553.390 108.020 ;
        RECT 616.010 107.820 616.330 107.880 ;
        RECT 2553.070 107.820 2553.390 107.880 ;
      LAYER via ;
        RECT 616.040 107.820 616.300 108.080 ;
        RECT 2553.100 107.820 2553.360 108.080 ;
      LAYER met2 ;
        RECT 615.830 500.000 616.110 504.000 ;
        RECT 615.870 498.850 616.010 500.000 ;
        RECT 615.870 498.710 616.240 498.850 ;
        RECT 616.100 108.110 616.240 498.710 ;
        RECT 616.040 107.790 616.300 108.110 ;
        RECT 2553.100 107.790 2553.360 108.110 ;
        RECT 2553.160 82.870 2553.300 107.790 ;
        RECT 2553.160 82.730 2555.600 82.870 ;
        RECT 2555.460 2.400 2555.600 82.730 ;
        RECT 2555.250 -4.800 2555.810 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.160 499.500 617.480 499.760 ;
        RECT 615.550 498.000 615.870 498.060 ;
        RECT 617.250 498.000 617.390 499.500 ;
        RECT 615.550 497.860 617.390 498.000 ;
        RECT 615.550 497.800 615.870 497.860 ;
        RECT 615.550 107.680 615.870 107.740 ;
        RECT 2566.870 107.680 2567.190 107.740 ;
        RECT 615.550 107.540 2567.190 107.680 ;
        RECT 615.550 107.480 615.870 107.540 ;
        RECT 2566.870 107.480 2567.190 107.540 ;
      LAYER via ;
        RECT 617.190 499.500 617.450 499.760 ;
        RECT 615.580 497.800 615.840 498.060 ;
        RECT 615.580 107.480 615.840 107.740 ;
        RECT 2566.900 107.480 2567.160 107.740 ;
      LAYER met2 ;
        RECT 617.210 500.000 617.490 504.000 ;
        RECT 617.250 499.790 617.390 500.000 ;
        RECT 617.190 499.470 617.450 499.790 ;
        RECT 615.580 497.770 615.840 498.090 ;
        RECT 615.640 107.770 615.780 497.770 ;
        RECT 615.580 107.450 615.840 107.770 ;
        RECT 2566.900 107.450 2567.160 107.770 ;
        RECT 2566.960 82.870 2567.100 107.450 ;
        RECT 2566.960 82.730 2572.160 82.870 ;
        RECT 2572.020 2.400 2572.160 82.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 618.540 499.160 618.860 499.420 ;
        RECT 616.930 497.320 617.250 497.380 ;
        RECT 618.630 497.320 618.770 499.160 ;
        RECT 616.930 497.180 618.770 497.320 ;
        RECT 616.930 497.120 617.250 497.180 ;
        RECT 614.630 472.160 614.950 472.220 ;
        RECT 616.470 472.160 616.790 472.220 ;
        RECT 614.630 472.020 616.790 472.160 ;
        RECT 614.630 471.960 614.950 472.020 ;
        RECT 616.470 471.960 616.790 472.020 ;
        RECT 614.630 31.860 614.950 31.920 ;
        RECT 2588.490 31.860 2588.810 31.920 ;
        RECT 614.630 31.720 2588.810 31.860 ;
        RECT 614.630 31.660 614.950 31.720 ;
        RECT 2588.490 31.660 2588.810 31.720 ;
      LAYER via ;
        RECT 618.570 499.160 618.830 499.420 ;
        RECT 616.960 497.120 617.220 497.380 ;
        RECT 614.660 471.960 614.920 472.220 ;
        RECT 616.500 471.960 616.760 472.220 ;
        RECT 614.660 31.660 614.920 31.920 ;
        RECT 2588.520 31.660 2588.780 31.920 ;
      LAYER met2 ;
        RECT 618.590 500.000 618.870 504.000 ;
        RECT 618.630 499.450 618.770 500.000 ;
        RECT 618.570 499.130 618.830 499.450 ;
        RECT 616.960 497.090 617.220 497.410 ;
        RECT 617.020 472.330 617.160 497.090 ;
        RECT 616.560 472.250 617.160 472.330 ;
        RECT 614.660 471.930 614.920 472.250 ;
        RECT 616.500 472.190 617.160 472.250 ;
        RECT 616.500 471.930 616.760 472.190 ;
        RECT 614.720 31.950 614.860 471.930 ;
        RECT 614.660 31.630 614.920 31.950 ;
        RECT 2588.520 31.630 2588.780 31.950 ;
        RECT 2588.580 2.400 2588.720 31.630 ;
        RECT 2588.370 -4.800 2588.930 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 619.920 499.500 620.240 499.760 ;
        RECT 620.010 499.020 620.150 499.500 ;
        RECT 619.780 498.880 620.150 499.020 ;
        RECT 619.780 498.400 619.920 498.880 ;
        RECT 619.690 498.140 620.010 498.400 ;
      LAYER via ;
        RECT 619.950 499.500 620.210 499.760 ;
        RECT 619.720 498.140 619.980 498.400 ;
      LAYER met2 ;
        RECT 619.970 500.000 620.250 504.000 ;
        RECT 620.010 499.790 620.150 500.000 ;
        RECT 619.950 499.470 620.210 499.790 ;
        RECT 619.720 498.110 619.980 498.430 ;
        RECT 619.780 488.085 619.920 498.110 ;
        RECT 619.710 487.715 619.990 488.085 ;
        RECT 2601.390 106.235 2601.670 106.605 ;
        RECT 2601.460 82.870 2601.600 106.235 ;
        RECT 2601.460 82.730 2605.280 82.870 ;
        RECT 2605.140 2.400 2605.280 82.730 ;
        RECT 2604.930 -4.800 2605.490 2.400 ;
      LAYER via2 ;
        RECT 619.710 487.760 619.990 488.040 ;
        RECT 2601.390 106.280 2601.670 106.560 ;
      LAYER met3 ;
        RECT 614.830 488.050 615.210 488.060 ;
        RECT 619.685 488.050 620.015 488.065 ;
        RECT 614.830 487.750 620.015 488.050 ;
        RECT 614.830 487.740 615.210 487.750 ;
        RECT 619.685 487.735 620.015 487.750 ;
        RECT 614.830 106.570 615.210 106.580 ;
        RECT 2601.365 106.570 2601.695 106.585 ;
        RECT 614.830 106.270 2601.695 106.570 ;
        RECT 614.830 106.260 615.210 106.270 ;
        RECT 2601.365 106.255 2601.695 106.270 ;
      LAYER via3 ;
        RECT 614.860 487.740 615.180 488.060 ;
        RECT 614.860 106.260 615.180 106.580 ;
      LAYER met4 ;
        RECT 614.855 487.735 615.185 488.065 ;
        RECT 614.870 106.585 615.170 487.735 ;
        RECT 614.855 106.255 615.185 106.585 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 471.480 622.310 471.540 ;
        RECT 623.830 471.480 624.150 471.540 ;
        RECT 621.990 471.340 624.150 471.480 ;
        RECT 621.990 471.280 622.310 471.340 ;
        RECT 623.830 471.280 624.150 471.340 ;
        RECT 623.830 107.340 624.150 107.400 ;
        RECT 2615.630 107.340 2615.950 107.400 ;
        RECT 623.830 107.200 2615.950 107.340 ;
        RECT 623.830 107.140 624.150 107.200 ;
        RECT 2615.630 107.140 2615.950 107.200 ;
        RECT 2615.630 37.640 2615.950 37.700 ;
        RECT 2621.610 37.640 2621.930 37.700 ;
        RECT 2615.630 37.500 2621.930 37.640 ;
        RECT 2615.630 37.440 2615.950 37.500 ;
        RECT 2621.610 37.440 2621.930 37.500 ;
      LAYER via ;
        RECT 622.020 471.280 622.280 471.540 ;
        RECT 623.860 471.280 624.120 471.540 ;
        RECT 623.860 107.140 624.120 107.400 ;
        RECT 2615.660 107.140 2615.920 107.400 ;
        RECT 2615.660 37.440 2615.920 37.700 ;
        RECT 2621.640 37.440 2621.900 37.700 ;
      LAYER met2 ;
        RECT 621.350 500.000 621.630 504.000 ;
        RECT 621.390 499.645 621.530 500.000 ;
        RECT 621.320 499.275 621.600 499.645 ;
        RECT 622.010 497.915 622.290 498.285 ;
        RECT 622.080 471.570 622.220 497.915 ;
        RECT 622.020 471.250 622.280 471.570 ;
        RECT 623.860 471.250 624.120 471.570 ;
        RECT 623.920 107.430 624.060 471.250 ;
        RECT 623.860 107.110 624.120 107.430 ;
        RECT 2615.660 107.110 2615.920 107.430 ;
        RECT 2615.720 37.730 2615.860 107.110 ;
        RECT 2615.660 37.410 2615.920 37.730 ;
        RECT 2621.640 37.410 2621.900 37.730 ;
        RECT 2621.700 2.400 2621.840 37.410 ;
        RECT 2621.490 -4.800 2622.050 2.400 ;
      LAYER via2 ;
        RECT 621.320 499.320 621.600 499.600 ;
        RECT 622.010 497.960 622.290 498.240 ;
      LAYER met3 ;
        RECT 621.295 499.295 621.625 499.625 ;
        RECT 621.310 498.250 621.610 499.295 ;
        RECT 621.985 498.250 622.315 498.265 ;
        RECT 621.310 497.950 622.315 498.250 ;
        RECT 621.985 497.935 622.315 497.950 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.910 38.660 623.230 38.720 ;
        RECT 2638.170 38.660 2638.490 38.720 ;
        RECT 622.910 38.520 2638.490 38.660 ;
        RECT 622.910 38.460 623.230 38.520 ;
        RECT 2638.170 38.460 2638.490 38.520 ;
      LAYER via ;
        RECT 622.940 38.460 623.200 38.720 ;
        RECT 2638.200 38.460 2638.460 38.720 ;
      LAYER met2 ;
        RECT 622.730 500.000 623.010 504.000 ;
        RECT 622.770 498.850 622.910 500.000 ;
        RECT 622.770 498.710 623.140 498.850 ;
        RECT 623.000 38.750 623.140 498.710 ;
        RECT 622.940 38.430 623.200 38.750 ;
        RECT 2638.200 38.430 2638.460 38.750 ;
        RECT 2638.260 2.400 2638.400 38.430 ;
        RECT 2638.050 -4.800 2638.610 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 472.160 622.770 472.220 ;
        RECT 623.830 472.160 624.150 472.220 ;
        RECT 622.450 472.020 624.150 472.160 ;
        RECT 622.450 471.960 622.770 472.020 ;
        RECT 623.830 471.960 624.150 472.020 ;
        RECT 622.450 38.320 622.770 38.380 ;
        RECT 2654.730 38.320 2655.050 38.380 ;
        RECT 622.450 38.180 2655.050 38.320 ;
        RECT 622.450 38.120 622.770 38.180 ;
        RECT 2654.730 38.120 2655.050 38.180 ;
      LAYER via ;
        RECT 622.480 471.960 622.740 472.220 ;
        RECT 623.860 471.960 624.120 472.220 ;
        RECT 622.480 38.120 622.740 38.380 ;
        RECT 2654.760 38.120 2655.020 38.380 ;
      LAYER met2 ;
        RECT 624.110 500.000 624.390 504.000 ;
        RECT 624.150 499.530 624.290 500.000 ;
        RECT 623.920 499.390 624.290 499.530 ;
        RECT 623.920 472.250 624.060 499.390 ;
        RECT 622.480 471.930 622.740 472.250 ;
        RECT 623.860 471.930 624.120 472.250 ;
        RECT 622.540 38.410 622.680 471.930 ;
        RECT 622.480 38.090 622.740 38.410 ;
        RECT 2654.760 38.090 2655.020 38.410 ;
        RECT 2654.820 2.400 2654.960 38.090 ;
        RECT 2654.610 -4.800 2655.170 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 470.800 622.310 470.860 ;
        RECT 625.210 470.800 625.530 470.860 ;
        RECT 621.990 470.660 625.530 470.800 ;
        RECT 621.990 470.600 622.310 470.660 ;
        RECT 625.210 470.600 625.530 470.660 ;
        RECT 621.990 37.980 622.310 38.040 ;
        RECT 2671.290 37.980 2671.610 38.040 ;
        RECT 621.990 37.840 2671.610 37.980 ;
        RECT 621.990 37.780 622.310 37.840 ;
        RECT 2671.290 37.780 2671.610 37.840 ;
      LAYER via ;
        RECT 622.020 470.600 622.280 470.860 ;
        RECT 625.240 470.600 625.500 470.860 ;
        RECT 622.020 37.780 622.280 38.040 ;
        RECT 2671.320 37.780 2671.580 38.040 ;
      LAYER met2 ;
        RECT 625.490 500.000 625.770 504.000 ;
        RECT 625.530 498.000 625.670 500.000 ;
        RECT 625.300 497.860 625.670 498.000 ;
        RECT 625.300 470.890 625.440 497.860 ;
        RECT 622.020 470.570 622.280 470.890 ;
        RECT 625.240 470.570 625.500 470.890 ;
        RECT 622.080 38.070 622.220 470.570 ;
        RECT 622.020 37.750 622.280 38.070 ;
        RECT 2671.320 37.750 2671.580 38.070 ;
        RECT 2671.380 2.400 2671.520 37.750 ;
        RECT 2671.170 -4.800 2671.730 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 492.560 476.490 492.620 ;
        RECT 477.090 492.560 477.410 492.620 ;
        RECT 476.170 492.420 477.410 492.560 ;
        RECT 476.170 492.360 476.490 492.420 ;
        RECT 477.090 492.360 477.410 492.420 ;
        RECT 477.090 109.040 477.410 109.100 ;
        RECT 876.830 109.040 877.150 109.100 ;
        RECT 477.090 108.900 877.150 109.040 ;
        RECT 477.090 108.840 477.410 108.900 ;
        RECT 876.830 108.840 877.150 108.900 ;
        RECT 876.830 20.300 877.150 20.360 ;
        RECT 882.810 20.300 883.130 20.360 ;
        RECT 876.830 20.160 883.130 20.300 ;
        RECT 876.830 20.100 877.150 20.160 ;
        RECT 882.810 20.100 883.130 20.160 ;
      LAYER via ;
        RECT 476.200 492.360 476.460 492.620 ;
        RECT 477.120 492.360 477.380 492.620 ;
        RECT 477.120 108.840 477.380 109.100 ;
        RECT 876.860 108.840 877.120 109.100 ;
        RECT 876.860 20.100 877.120 20.360 ;
        RECT 882.840 20.100 883.100 20.360 ;
      LAYER met2 ;
        RECT 476.450 500.000 476.730 504.000 ;
        RECT 476.490 498.340 476.630 500.000 ;
        RECT 476.260 498.200 476.630 498.340 ;
        RECT 476.260 492.650 476.400 498.200 ;
        RECT 476.200 492.330 476.460 492.650 ;
        RECT 477.120 492.330 477.380 492.650 ;
        RECT 477.180 109.130 477.320 492.330 ;
        RECT 477.120 108.810 477.380 109.130 ;
        RECT 876.860 108.810 877.120 109.130 ;
        RECT 876.920 20.390 877.060 108.810 ;
        RECT 876.860 20.070 877.120 20.390 ;
        RECT 882.840 20.070 883.100 20.390 ;
        RECT 882.900 2.400 883.040 20.070 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.870 500.000 627.150 504.000 ;
        RECT 626.910 498.850 627.050 500.000 ;
        RECT 626.680 498.710 627.050 498.850 ;
        RECT 626.680 483.325 626.820 498.710 ;
        RECT 626.610 482.955 626.890 483.325 ;
        RECT 2684.190 113.715 2684.470 114.085 ;
        RECT 2684.260 82.870 2684.400 113.715 ;
        RECT 2684.260 82.730 2688.080 82.870 ;
        RECT 2687.940 2.400 2688.080 82.730 ;
        RECT 2687.730 -4.800 2688.290 2.400 ;
      LAYER via2 ;
        RECT 626.610 483.000 626.890 483.280 ;
        RECT 2684.190 113.760 2684.470 114.040 ;
      LAYER met3 ;
        RECT 625.870 483.290 626.250 483.300 ;
        RECT 626.585 483.290 626.915 483.305 ;
        RECT 625.870 482.990 626.915 483.290 ;
        RECT 625.870 482.980 626.250 482.990 ;
        RECT 626.585 482.975 626.915 482.990 ;
        RECT 625.870 114.050 626.250 114.060 ;
        RECT 2684.165 114.050 2684.495 114.065 ;
        RECT 625.870 113.750 2684.495 114.050 ;
        RECT 625.870 113.740 626.250 113.750 ;
        RECT 2684.165 113.735 2684.495 113.750 ;
      LAYER via3 ;
        RECT 625.900 482.980 626.220 483.300 ;
        RECT 625.900 113.740 626.220 114.060 ;
      LAYER met4 ;
        RECT 625.895 482.975 626.225 483.305 ;
        RECT 625.910 114.065 626.210 482.975 ;
        RECT 625.895 113.735 626.225 114.065 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.890 51.580 629.210 51.640 ;
        RECT 2697.970 51.580 2698.290 51.640 ;
        RECT 628.890 51.440 2698.290 51.580 ;
        RECT 628.890 51.380 629.210 51.440 ;
        RECT 2697.970 51.380 2698.290 51.440 ;
        RECT 2697.970 17.580 2698.290 17.640 ;
        RECT 2704.410 17.580 2704.730 17.640 ;
        RECT 2697.970 17.440 2704.730 17.580 ;
        RECT 2697.970 17.380 2698.290 17.440 ;
        RECT 2704.410 17.380 2704.730 17.440 ;
      LAYER via ;
        RECT 628.920 51.380 629.180 51.640 ;
        RECT 2698.000 51.380 2698.260 51.640 ;
        RECT 2698.000 17.380 2698.260 17.640 ;
        RECT 2704.440 17.380 2704.700 17.640 ;
      LAYER met2 ;
        RECT 628.250 500.000 628.530 504.000 ;
        RECT 628.290 499.815 628.430 500.000 ;
        RECT 628.220 499.445 628.500 499.815 ;
        RECT 628.910 497.235 629.190 497.605 ;
        RECT 628.980 51.670 629.120 497.235 ;
        RECT 628.920 51.350 629.180 51.670 ;
        RECT 2698.000 51.350 2698.260 51.670 ;
        RECT 2698.060 17.670 2698.200 51.350 ;
        RECT 2698.000 17.350 2698.260 17.670 ;
        RECT 2704.440 17.350 2704.700 17.670 ;
        RECT 2704.500 2.400 2704.640 17.350 ;
        RECT 2704.290 -4.800 2704.850 2.400 ;
      LAYER via2 ;
        RECT 628.220 499.490 628.500 499.770 ;
        RECT 628.910 497.280 629.190 497.560 ;
      LAYER met3 ;
        RECT 628.195 499.465 628.525 499.795 ;
        RECT 628.210 497.570 628.510 499.465 ;
        RECT 628.885 497.570 629.215 497.585 ;
        RECT 628.210 497.270 629.215 497.570 ;
        RECT 628.885 497.255 629.215 497.270 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.350 58.720 629.670 58.780 ;
        RECT 2720.970 58.720 2721.290 58.780 ;
        RECT 629.350 58.580 2721.290 58.720 ;
        RECT 629.350 58.520 629.670 58.580 ;
        RECT 2720.970 58.520 2721.290 58.580 ;
      LAYER via ;
        RECT 629.380 58.520 629.640 58.780 ;
        RECT 2721.000 58.520 2721.260 58.780 ;
      LAYER met2 ;
        RECT 629.630 500.000 629.910 504.000 ;
        RECT 629.670 499.815 629.810 500.000 ;
        RECT 629.600 499.445 629.880 499.815 ;
        RECT 629.370 497.915 629.650 498.285 ;
        RECT 629.440 58.810 629.580 497.915 ;
        RECT 629.380 58.490 629.640 58.810 ;
        RECT 2721.000 58.490 2721.260 58.810 ;
        RECT 2721.060 2.400 2721.200 58.490 ;
        RECT 2720.850 -4.800 2721.410 2.400 ;
      LAYER via2 ;
        RECT 629.600 499.490 629.880 499.770 ;
        RECT 629.370 497.960 629.650 498.240 ;
      LAYER met3 ;
        RECT 629.575 499.465 629.905 499.795 ;
        RECT 629.590 498.265 629.890 499.465 ;
        RECT 629.345 497.950 629.890 498.265 ;
        RECT 629.345 497.935 629.675 497.950 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.270 100.540 630.590 100.600 ;
        RECT 2732.470 100.540 2732.790 100.600 ;
        RECT 630.270 100.400 2732.790 100.540 ;
        RECT 630.270 100.340 630.590 100.400 ;
        RECT 2732.470 100.340 2732.790 100.400 ;
      LAYER via ;
        RECT 630.300 100.340 630.560 100.600 ;
        RECT 2732.500 100.340 2732.760 100.600 ;
      LAYER met2 ;
        RECT 631.010 500.000 631.290 504.000 ;
        RECT 631.050 499.815 631.190 500.000 ;
        RECT 630.980 499.445 631.260 499.815 ;
        RECT 630.290 491.115 630.570 491.485 ;
        RECT 630.360 100.630 630.500 491.115 ;
        RECT 630.300 100.310 630.560 100.630 ;
        RECT 2732.500 100.310 2732.760 100.630 ;
        RECT 2732.560 82.870 2732.700 100.310 ;
        RECT 2732.560 82.730 2737.760 82.870 ;
        RECT 2737.620 2.400 2737.760 82.730 ;
        RECT 2737.410 -4.800 2737.970 2.400 ;
      LAYER via2 ;
        RECT 630.980 499.490 631.260 499.770 ;
        RECT 630.290 491.160 630.570 491.440 ;
      LAYER met3 ;
        RECT 630.955 499.780 631.285 499.795 ;
        RECT 630.740 499.620 631.285 499.780 ;
        RECT 630.470 499.465 631.285 499.620 ;
        RECT 630.470 499.310 631.040 499.465 ;
        RECT 630.470 499.300 630.850 499.310 ;
        RECT 630.265 491.460 630.595 491.465 ;
        RECT 630.265 491.450 630.850 491.460 ;
        RECT 630.040 491.150 630.850 491.450 ;
        RECT 630.265 491.140 630.850 491.150 ;
        RECT 630.265 491.135 630.595 491.140 ;
      LAYER via3 ;
        RECT 630.500 499.300 630.820 499.620 ;
        RECT 630.500 491.140 630.820 491.460 ;
      LAYER met4 ;
        RECT 630.495 499.295 630.825 499.625 ;
        RECT 630.510 491.465 630.810 499.295 ;
        RECT 630.495 491.135 630.825 491.465 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.730 107.000 631.050 107.060 ;
        RECT 2753.170 107.000 2753.490 107.060 ;
        RECT 630.730 106.860 2753.490 107.000 ;
        RECT 630.730 106.800 631.050 106.860 ;
        RECT 2753.170 106.800 2753.490 106.860 ;
      LAYER via ;
        RECT 630.760 106.800 631.020 107.060 ;
        RECT 2753.200 106.800 2753.460 107.060 ;
      LAYER met2 ;
        RECT 632.390 500.000 632.670 504.000 ;
        RECT 632.430 499.815 632.570 500.000 ;
        RECT 632.360 499.445 632.640 499.815 ;
        RECT 630.750 495.875 631.030 496.245 ;
        RECT 630.820 107.090 630.960 495.875 ;
        RECT 630.760 106.770 631.020 107.090 ;
        RECT 2753.200 106.770 2753.460 107.090 ;
        RECT 2753.260 17.410 2753.400 106.770 ;
        RECT 2753.260 17.270 2754.320 17.410 ;
        RECT 2754.180 2.400 2754.320 17.270 ;
        RECT 2753.970 -4.800 2754.530 2.400 ;
      LAYER via2 ;
        RECT 632.360 499.490 632.640 499.770 ;
        RECT 630.750 495.920 631.030 496.200 ;
      LAYER met3 ;
        RECT 632.335 499.465 632.665 499.795 ;
        RECT 630.725 496.210 631.055 496.225 ;
        RECT 632.350 496.210 632.650 499.465 ;
        RECT 630.725 495.910 632.650 496.210 ;
        RECT 630.725 495.895 631.055 495.910 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.770 500.000 634.050 504.000 ;
        RECT 633.810 498.340 633.950 500.000 ;
        RECT 633.580 498.200 633.950 498.340 ;
        RECT 633.580 490.805 633.720 498.200 ;
        RECT 633.510 490.435 633.790 490.805 ;
        RECT 2766.990 113.035 2767.270 113.405 ;
        RECT 2767.060 82.870 2767.200 113.035 ;
        RECT 2767.060 82.730 2770.880 82.870 ;
        RECT 2770.740 2.400 2770.880 82.730 ;
        RECT 2770.530 -4.800 2771.090 2.400 ;
      LAYER via2 ;
        RECT 633.510 490.480 633.790 490.760 ;
        RECT 2766.990 113.080 2767.270 113.360 ;
      LAYER met3 ;
        RECT 633.485 490.780 633.815 490.785 ;
        RECT 633.230 490.770 633.815 490.780 ;
        RECT 633.030 490.470 633.815 490.770 ;
        RECT 633.230 490.460 633.815 490.470 ;
        RECT 633.485 490.455 633.815 490.460 ;
        RECT 633.230 113.370 633.610 113.380 ;
        RECT 2766.965 113.370 2767.295 113.385 ;
        RECT 633.230 113.070 2767.295 113.370 ;
        RECT 633.230 113.060 633.610 113.070 ;
        RECT 2766.965 113.055 2767.295 113.070 ;
      LAYER via3 ;
        RECT 633.260 490.460 633.580 490.780 ;
        RECT 633.260 113.060 633.580 113.380 ;
      LAYER met4 ;
        RECT 633.255 490.455 633.585 490.785 ;
        RECT 633.270 113.385 633.570 490.455 ;
        RECT 633.255 113.055 633.585 113.385 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.100 499.500 635.420 499.760 ;
        RECT 635.190 498.740 635.330 499.500 ;
        RECT 635.190 498.540 635.650 498.740 ;
        RECT 635.330 498.480 635.650 498.540 ;
        RECT 635.330 487.460 635.650 487.520 ;
        RECT 1045.190 487.460 1045.510 487.520 ;
        RECT 635.330 487.320 1045.510 487.460 ;
        RECT 635.330 487.260 635.650 487.320 ;
        RECT 1045.190 487.260 1045.510 487.320 ;
        RECT 1045.190 44.780 1045.510 44.840 ;
        RECT 2787.210 44.780 2787.530 44.840 ;
        RECT 1045.190 44.640 2787.530 44.780 ;
        RECT 1045.190 44.580 1045.510 44.640 ;
        RECT 2787.210 44.580 2787.530 44.640 ;
      LAYER via ;
        RECT 635.130 499.500 635.390 499.760 ;
        RECT 635.360 498.480 635.620 498.740 ;
        RECT 635.360 487.260 635.620 487.520 ;
        RECT 1045.220 487.260 1045.480 487.520 ;
        RECT 1045.220 44.580 1045.480 44.840 ;
        RECT 2787.240 44.580 2787.500 44.840 ;
      LAYER met2 ;
        RECT 635.150 500.000 635.430 504.000 ;
        RECT 635.190 499.790 635.330 500.000 ;
        RECT 635.130 499.470 635.390 499.790 ;
        RECT 635.360 498.450 635.620 498.770 ;
        RECT 635.420 487.550 635.560 498.450 ;
        RECT 635.360 487.230 635.620 487.550 ;
        RECT 1045.220 487.230 1045.480 487.550 ;
        RECT 1045.280 44.870 1045.420 487.230 ;
        RECT 1045.220 44.550 1045.480 44.870 ;
        RECT 2787.240 44.550 2787.500 44.870 ;
        RECT 2787.300 2.400 2787.440 44.550 ;
        RECT 2787.090 -4.800 2787.650 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.710 491.540 637.030 491.600 ;
        RECT 638.550 491.540 638.870 491.600 ;
        RECT 636.710 491.400 638.870 491.540 ;
        RECT 636.710 491.340 637.030 491.400 ;
        RECT 638.550 491.340 638.870 491.400 ;
        RECT 638.550 79.460 638.870 79.520 ;
        RECT 2803.770 79.460 2804.090 79.520 ;
        RECT 638.550 79.320 2804.090 79.460 ;
        RECT 638.550 79.260 638.870 79.320 ;
        RECT 2803.770 79.260 2804.090 79.320 ;
      LAYER via ;
        RECT 636.740 491.340 637.000 491.600 ;
        RECT 638.580 491.340 638.840 491.600 ;
        RECT 638.580 79.260 638.840 79.520 ;
        RECT 2803.800 79.260 2804.060 79.520 ;
      LAYER met2 ;
        RECT 636.530 500.000 636.810 504.000 ;
        RECT 636.570 498.680 636.710 500.000 ;
        RECT 636.570 498.540 636.940 498.680 ;
        RECT 636.800 491.630 636.940 498.540 ;
        RECT 636.740 491.310 637.000 491.630 ;
        RECT 638.580 491.310 638.840 491.630 ;
        RECT 638.640 79.550 638.780 491.310 ;
        RECT 638.580 79.230 638.840 79.550 ;
        RECT 2803.800 79.230 2804.060 79.550 ;
        RECT 2803.860 2.400 2804.000 79.230 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.010 115.840 478.330 115.900 ;
        RECT 897.070 115.840 897.390 115.900 ;
        RECT 478.010 115.700 897.390 115.840 ;
        RECT 478.010 115.640 478.330 115.700 ;
        RECT 897.070 115.640 897.390 115.700 ;
      LAYER via ;
        RECT 478.040 115.640 478.300 115.900 ;
        RECT 897.100 115.640 897.360 115.900 ;
      LAYER met2 ;
        RECT 477.830 500.000 478.110 504.000 ;
        RECT 477.870 499.020 478.010 500.000 ;
        RECT 477.640 498.880 478.010 499.020 ;
        RECT 477.640 498.340 477.780 498.880 ;
        RECT 477.640 498.200 478.240 498.340 ;
        RECT 478.100 115.930 478.240 498.200 ;
        RECT 478.040 115.610 478.300 115.930 ;
        RECT 897.100 115.610 897.360 115.930 ;
        RECT 897.160 82.870 897.300 115.610 ;
        RECT 897.160 82.730 899.600 82.870 ;
        RECT 899.460 2.400 899.600 82.730 ;
        RECT 899.250 -4.800 899.810 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.550 472.840 477.870 472.900 ;
        RECT 478.930 472.840 479.250 472.900 ;
        RECT 477.550 472.700 479.250 472.840 ;
        RECT 477.550 472.640 477.870 472.700 ;
        RECT 478.930 472.640 479.250 472.700 ;
        RECT 477.550 115.500 477.870 115.560 ;
        RECT 910.870 115.500 911.190 115.560 ;
        RECT 477.550 115.360 911.190 115.500 ;
        RECT 477.550 115.300 477.870 115.360 ;
        RECT 910.870 115.300 911.190 115.360 ;
      LAYER via ;
        RECT 477.580 472.640 477.840 472.900 ;
        RECT 478.960 472.640 479.220 472.900 ;
        RECT 477.580 115.300 477.840 115.560 ;
        RECT 910.900 115.300 911.160 115.560 ;
      LAYER met2 ;
        RECT 479.210 500.000 479.490 504.000 ;
        RECT 479.250 498.850 479.390 500.000 ;
        RECT 479.020 498.710 479.390 498.850 ;
        RECT 479.020 472.930 479.160 498.710 ;
        RECT 477.580 472.610 477.840 472.930 ;
        RECT 478.960 472.610 479.220 472.930 ;
        RECT 477.640 115.590 477.780 472.610 ;
        RECT 477.580 115.270 477.840 115.590 ;
        RECT 910.900 115.270 911.160 115.590 ;
        RECT 910.960 82.870 911.100 115.270 ;
        RECT 910.960 82.730 916.160 82.870 ;
        RECT 916.020 2.400 916.160 82.730 ;
        RECT 915.810 -4.800 916.370 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 481.230 27.100 481.550 27.160 ;
        RECT 481.230 26.960 517.570 27.100 ;
        RECT 481.230 26.900 481.550 26.960 ;
        RECT 517.430 26.760 517.570 26.960 ;
        RECT 932.490 26.760 932.810 26.820 ;
        RECT 517.430 26.620 932.810 26.760 ;
        RECT 932.490 26.560 932.810 26.620 ;
      LAYER via ;
        RECT 481.260 26.900 481.520 27.160 ;
        RECT 932.520 26.560 932.780 26.820 ;
      LAYER met2 ;
        RECT 480.590 500.000 480.870 504.000 ;
        RECT 480.630 498.680 480.770 500.000 ;
        RECT 480.630 498.540 481.460 498.680 ;
        RECT 481.320 27.190 481.460 498.540 ;
        RECT 481.260 26.870 481.520 27.190 ;
        RECT 932.520 26.530 932.780 26.850 ;
        RECT 932.580 2.400 932.720 26.530 ;
        RECT 932.370 -4.800 932.930 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.970 500.000 482.250 504.000 ;
        RECT 482.010 498.965 482.150 500.000 ;
        RECT 481.940 498.595 482.220 498.965 ;
        RECT 949.070 37.555 949.350 37.925 ;
        RECT 949.140 2.400 949.280 37.555 ;
        RECT 948.930 -4.800 949.490 2.400 ;
      LAYER via2 ;
        RECT 481.940 498.640 482.220 498.920 ;
        RECT 949.070 37.600 949.350 37.880 ;
      LAYER met3 ;
        RECT 480.510 498.930 480.890 498.940 ;
        RECT 481.915 498.930 482.245 498.945 ;
        RECT 480.510 498.630 482.245 498.930 ;
        RECT 480.510 498.620 480.890 498.630 ;
        RECT 481.915 498.615 482.245 498.630 ;
        RECT 480.510 37.890 480.890 37.900 ;
        RECT 949.045 37.890 949.375 37.905 ;
        RECT 480.510 37.590 949.375 37.890 ;
        RECT 480.510 37.580 480.890 37.590 ;
        RECT 949.045 37.575 949.375 37.590 ;
      LAYER via3 ;
        RECT 480.540 498.620 480.860 498.940 ;
        RECT 480.540 37.580 480.860 37.900 ;
      LAYER met4 ;
        RECT 480.535 498.615 480.865 498.945 ;
        RECT 480.550 37.905 480.850 498.615 ;
        RECT 480.535 37.575 480.865 37.905 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.990 473.320 484.310 473.580 ;
        RECT 484.080 472.560 484.220 473.320 ;
        RECT 483.990 472.300 484.310 472.560 ;
        RECT 483.990 115.160 484.310 115.220 ;
        RECT 959.630 115.160 959.950 115.220 ;
        RECT 483.990 115.020 959.950 115.160 ;
        RECT 483.990 114.960 484.310 115.020 ;
        RECT 959.630 114.960 959.950 115.020 ;
        RECT 959.630 20.300 959.950 20.360 ;
        RECT 965.610 20.300 965.930 20.360 ;
        RECT 959.630 20.160 965.930 20.300 ;
        RECT 959.630 20.100 959.950 20.160 ;
        RECT 965.610 20.100 965.930 20.160 ;
      LAYER via ;
        RECT 484.020 473.320 484.280 473.580 ;
        RECT 484.020 472.300 484.280 472.560 ;
        RECT 484.020 114.960 484.280 115.220 ;
        RECT 959.660 114.960 959.920 115.220 ;
        RECT 959.660 20.100 959.920 20.360 ;
        RECT 965.640 20.100 965.900 20.360 ;
      LAYER met2 ;
        RECT 483.350 500.000 483.630 504.000 ;
        RECT 483.390 499.020 483.530 500.000 ;
        RECT 483.390 498.880 483.990 499.020 ;
        RECT 483.850 498.850 483.990 498.880 ;
        RECT 483.850 498.710 484.220 498.850 ;
        RECT 484.080 473.610 484.220 498.710 ;
        RECT 484.020 473.290 484.280 473.610 ;
        RECT 484.020 472.270 484.280 472.590 ;
        RECT 484.080 115.250 484.220 472.270 ;
        RECT 484.020 114.930 484.280 115.250 ;
        RECT 959.660 114.930 959.920 115.250 ;
        RECT 959.720 20.390 959.860 114.930 ;
        RECT 959.660 20.070 959.920 20.390 ;
        RECT 965.640 20.070 965.900 20.390 ;
        RECT 965.700 2.400 965.840 20.070 ;
        RECT 965.490 -4.800 966.050 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.680 499.500 485.000 499.760 ;
        RECT 484.770 498.740 484.910 499.500 ;
        RECT 484.450 498.540 484.910 498.740 ;
        RECT 484.450 498.480 484.770 498.540 ;
        RECT 483.530 114.820 483.850 114.880 ;
        RECT 979.870 114.820 980.190 114.880 ;
        RECT 483.530 114.680 980.190 114.820 ;
        RECT 483.530 114.620 483.850 114.680 ;
        RECT 979.870 114.620 980.190 114.680 ;
      LAYER via ;
        RECT 484.710 499.500 484.970 499.760 ;
        RECT 484.480 498.480 484.740 498.740 ;
        RECT 483.560 114.620 483.820 114.880 ;
        RECT 979.900 114.620 980.160 114.880 ;
      LAYER met2 ;
        RECT 484.730 500.000 485.010 504.000 ;
        RECT 484.770 499.790 484.910 500.000 ;
        RECT 484.710 499.470 484.970 499.790 ;
        RECT 484.480 498.450 484.740 498.770 ;
        RECT 484.540 473.010 484.680 498.450 ;
        RECT 483.620 472.870 484.680 473.010 ;
        RECT 483.620 114.910 483.760 472.870 ;
        RECT 483.560 114.590 483.820 114.910 ;
        RECT 979.900 114.590 980.160 114.910 ;
        RECT 979.960 82.870 980.100 114.590 ;
        RECT 979.960 82.730 982.400 82.870 ;
        RECT 982.260 2.400 982.400 82.730 ;
        RECT 982.050 -4.800 982.610 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.450 472.500 484.770 472.560 ;
        RECT 486.750 472.500 487.070 472.560 ;
        RECT 484.450 472.360 487.070 472.500 ;
        RECT 484.450 472.300 484.770 472.360 ;
        RECT 486.750 472.300 487.070 472.360 ;
        RECT 484.450 122.300 484.770 122.360 ;
        RECT 993.670 122.300 993.990 122.360 ;
        RECT 484.450 122.160 993.990 122.300 ;
        RECT 484.450 122.100 484.770 122.160 ;
        RECT 993.670 122.100 993.990 122.160 ;
      LAYER via ;
        RECT 484.480 472.300 484.740 472.560 ;
        RECT 486.780 472.300 487.040 472.560 ;
        RECT 484.480 122.100 484.740 122.360 ;
        RECT 993.700 122.100 993.960 122.360 ;
      LAYER met2 ;
        RECT 486.110 500.000 486.390 504.000 ;
        RECT 486.150 499.815 486.290 500.000 ;
        RECT 486.080 499.445 486.360 499.815 ;
        RECT 486.770 497.915 487.050 498.285 ;
        RECT 486.840 472.590 486.980 497.915 ;
        RECT 484.480 472.270 484.740 472.590 ;
        RECT 486.780 472.270 487.040 472.590 ;
        RECT 484.540 122.390 484.680 472.270 ;
        RECT 484.480 122.070 484.740 122.390 ;
        RECT 993.700 122.070 993.960 122.390 ;
        RECT 993.760 82.870 993.900 122.070 ;
        RECT 993.760 82.730 998.960 82.870 ;
        RECT 998.820 2.400 998.960 82.730 ;
        RECT 998.610 -4.800 999.170 2.400 ;
      LAYER via2 ;
        RECT 486.080 499.490 486.360 499.770 ;
        RECT 486.770 497.960 487.050 498.240 ;
      LAYER met3 ;
        RECT 486.055 499.465 486.385 499.795 ;
        RECT 486.070 498.250 486.370 499.465 ;
        RECT 486.745 498.250 487.075 498.265 ;
        RECT 486.070 497.950 487.075 498.250 ;
        RECT 486.745 497.935 487.075 497.950 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.490 500.000 487.770 504.000 ;
        RECT 487.530 499.700 487.670 500.000 ;
        RECT 487.530 499.560 487.900 499.700 ;
        RECT 487.760 498.965 487.900 499.560 ;
        RECT 487.690 498.595 487.970 498.965 ;
        RECT 1015.310 47.075 1015.590 47.445 ;
        RECT 1015.380 2.400 1015.520 47.075 ;
        RECT 1015.170 -4.800 1015.730 2.400 ;
      LAYER via2 ;
        RECT 487.690 498.640 487.970 498.920 ;
        RECT 1015.310 47.120 1015.590 47.400 ;
      LAYER met3 ;
        RECT 487.665 498.930 487.995 498.945 ;
        RECT 488.790 498.930 489.170 498.940 ;
        RECT 487.665 498.630 489.170 498.930 ;
        RECT 487.665 498.615 487.995 498.630 ;
        RECT 488.790 498.620 489.170 498.630 ;
        RECT 488.790 47.410 489.170 47.420 ;
        RECT 1015.285 47.410 1015.615 47.425 ;
        RECT 488.790 47.110 1015.615 47.410 ;
        RECT 488.790 47.100 489.170 47.110 ;
        RECT 1015.285 47.095 1015.615 47.110 ;
      LAYER via3 ;
        RECT 488.820 498.620 489.140 498.940 ;
        RECT 488.820 47.100 489.140 47.420 ;
      LAYER met4 ;
        RECT 488.815 498.615 489.145 498.945 ;
        RECT 488.830 47.425 489.130 498.615 ;
        RECT 488.815 47.095 489.145 47.425 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 122.640 463.610 122.700 ;
        RECT 711.230 122.640 711.550 122.700 ;
        RECT 463.290 122.500 711.550 122.640 ;
        RECT 463.290 122.440 463.610 122.500 ;
        RECT 711.230 122.440 711.550 122.500 ;
        RECT 711.230 19.960 711.550 20.020 ;
        RECT 717.210 19.960 717.530 20.020 ;
        RECT 711.230 19.820 717.530 19.960 ;
        RECT 711.230 19.760 711.550 19.820 ;
        RECT 717.210 19.760 717.530 19.820 ;
      LAYER via ;
        RECT 463.320 122.440 463.580 122.700 ;
        RECT 711.260 122.440 711.520 122.700 ;
        RECT 711.260 19.760 711.520 20.020 ;
        RECT 717.240 19.760 717.500 20.020 ;
      LAYER met2 ;
        RECT 462.650 500.000 462.930 504.000 ;
        RECT 462.690 498.680 462.830 500.000 ;
        RECT 462.690 498.540 463.520 498.680 ;
        RECT 463.380 122.730 463.520 498.540 ;
        RECT 463.320 122.410 463.580 122.730 ;
        RECT 711.260 122.410 711.520 122.730 ;
        RECT 711.320 20.050 711.460 122.410 ;
        RECT 711.260 19.730 711.520 20.050 ;
        RECT 717.240 19.730 717.500 20.050 ;
        RECT 717.300 2.400 717.440 19.730 ;
        RECT 717.090 -4.800 717.650 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 488.820 499.160 489.140 499.420 ;
        RECT 487.670 498.000 487.990 498.060 ;
        RECT 488.910 498.000 489.050 499.160 ;
        RECT 487.670 497.860 489.050 498.000 ;
        RECT 487.670 497.800 487.990 497.860 ;
      LAYER via ;
        RECT 488.850 499.160 489.110 499.420 ;
        RECT 487.700 497.800 487.960 498.060 ;
      LAYER met2 ;
        RECT 488.870 500.000 489.150 504.000 ;
        RECT 488.910 499.450 489.050 500.000 ;
        RECT 488.850 499.130 489.110 499.450 ;
        RECT 487.700 497.770 487.960 498.090 ;
        RECT 487.760 488.085 487.900 497.770 ;
        RECT 487.690 487.715 487.970 488.085 ;
        RECT 1031.870 46.395 1032.150 46.765 ;
        RECT 1031.940 2.400 1032.080 46.395 ;
        RECT 1031.730 -4.800 1032.290 2.400 ;
      LAYER via2 ;
        RECT 487.690 487.760 487.970 488.040 ;
        RECT 1031.870 46.440 1032.150 46.720 ;
      LAYER met3 ;
        RECT 487.665 488.060 487.995 488.065 ;
        RECT 487.665 488.050 488.250 488.060 ;
        RECT 487.665 487.750 488.450 488.050 ;
        RECT 487.665 487.740 488.250 487.750 ;
        RECT 487.665 487.735 487.995 487.740 ;
        RECT 487.870 46.730 488.250 46.740 ;
        RECT 1031.845 46.730 1032.175 46.745 ;
        RECT 487.870 46.430 1032.175 46.730 ;
        RECT 487.870 46.420 488.250 46.430 ;
        RECT 1031.845 46.415 1032.175 46.430 ;
      LAYER via3 ;
        RECT 487.900 487.740 488.220 488.060 ;
        RECT 487.900 46.420 488.220 46.740 ;
      LAYER met4 ;
        RECT 487.895 487.735 488.225 488.065 ;
        RECT 487.910 46.745 488.210 487.735 ;
        RECT 487.895 46.415 488.225 46.745 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.890 121.960 491.210 122.020 ;
        RECT 1042.430 121.960 1042.750 122.020 ;
        RECT 490.890 121.820 1042.750 121.960 ;
        RECT 490.890 121.760 491.210 121.820 ;
        RECT 1042.430 121.760 1042.750 121.820 ;
        RECT 1042.430 20.300 1042.750 20.360 ;
        RECT 1048.410 20.300 1048.730 20.360 ;
        RECT 1042.430 20.160 1048.730 20.300 ;
        RECT 1042.430 20.100 1042.750 20.160 ;
        RECT 1048.410 20.100 1048.730 20.160 ;
      LAYER via ;
        RECT 490.920 121.760 491.180 122.020 ;
        RECT 1042.460 121.760 1042.720 122.020 ;
        RECT 1042.460 20.100 1042.720 20.360 ;
        RECT 1048.440 20.100 1048.700 20.360 ;
      LAYER met2 ;
        RECT 490.250 500.000 490.530 504.000 ;
        RECT 490.290 499.815 490.430 500.000 ;
        RECT 490.220 499.445 490.500 499.815 ;
        RECT 490.910 487.715 491.190 488.085 ;
        RECT 490.980 122.050 491.120 487.715 ;
        RECT 490.920 121.730 491.180 122.050 ;
        RECT 1042.460 121.730 1042.720 122.050 ;
        RECT 1042.520 20.390 1042.660 121.730 ;
        RECT 1042.460 20.070 1042.720 20.390 ;
        RECT 1048.440 20.070 1048.700 20.390 ;
        RECT 1048.500 2.400 1048.640 20.070 ;
        RECT 1048.290 -4.800 1048.850 2.400 ;
      LAYER via2 ;
        RECT 490.220 499.490 490.500 499.770 ;
        RECT 490.910 487.760 491.190 488.040 ;
      LAYER met3 ;
        RECT 490.195 499.780 490.525 499.795 ;
        RECT 490.195 499.620 490.740 499.780 ;
        RECT 490.195 499.465 491.010 499.620 ;
        RECT 490.440 499.310 491.010 499.465 ;
        RECT 490.630 499.300 491.010 499.310 ;
        RECT 490.885 488.060 491.215 488.065 ;
        RECT 490.630 488.050 491.215 488.060 ;
        RECT 490.630 487.750 491.440 488.050 ;
        RECT 490.630 487.740 491.215 487.750 ;
        RECT 490.885 487.735 491.215 487.740 ;
      LAYER via3 ;
        RECT 490.660 499.300 490.980 499.620 ;
        RECT 490.660 487.740 490.980 488.060 ;
      LAYER met4 ;
        RECT 490.655 499.295 490.985 499.625 ;
        RECT 490.670 488.065 490.970 499.295 ;
        RECT 490.655 487.735 490.985 488.065 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 472.840 490.750 472.900 ;
        RECT 491.350 472.840 491.670 472.900 ;
        RECT 490.430 472.700 491.670 472.840 ;
        RECT 490.430 472.640 490.750 472.700 ;
        RECT 491.350 472.640 491.670 472.700 ;
        RECT 490.430 121.620 490.750 121.680 ;
        RECT 1062.670 121.620 1062.990 121.680 ;
        RECT 490.430 121.480 1062.990 121.620 ;
        RECT 490.430 121.420 490.750 121.480 ;
        RECT 1062.670 121.420 1062.990 121.480 ;
      LAYER via ;
        RECT 490.460 472.640 490.720 472.900 ;
        RECT 491.380 472.640 491.640 472.900 ;
        RECT 490.460 121.420 490.720 121.680 ;
        RECT 1062.700 121.420 1062.960 121.680 ;
      LAYER met2 ;
        RECT 491.630 500.000 491.910 504.000 ;
        RECT 491.670 499.815 491.810 500.000 ;
        RECT 491.600 499.445 491.880 499.815 ;
        RECT 491.370 497.915 491.650 498.285 ;
        RECT 491.440 472.930 491.580 497.915 ;
        RECT 490.460 472.610 490.720 472.930 ;
        RECT 491.380 472.610 491.640 472.930 ;
        RECT 490.520 121.710 490.660 472.610 ;
        RECT 490.460 121.390 490.720 121.710 ;
        RECT 1062.700 121.390 1062.960 121.710 ;
        RECT 1062.760 82.870 1062.900 121.390 ;
        RECT 1062.760 82.730 1065.200 82.870 ;
        RECT 1065.060 2.400 1065.200 82.730 ;
        RECT 1064.850 -4.800 1065.410 2.400 ;
      LAYER via2 ;
        RECT 491.600 499.490 491.880 499.770 ;
        RECT 491.370 497.960 491.650 498.240 ;
      LAYER met3 ;
        RECT 491.575 499.465 491.905 499.795 ;
        RECT 491.590 498.265 491.890 499.465 ;
        RECT 491.345 497.950 491.890 498.265 ;
        RECT 491.345 497.935 491.675 497.950 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 491.350 121.280 491.670 121.340 ;
        RECT 1076.470 121.280 1076.790 121.340 ;
        RECT 491.350 121.140 1076.790 121.280 ;
        RECT 491.350 121.080 491.670 121.140 ;
        RECT 1076.470 121.080 1076.790 121.140 ;
      LAYER via ;
        RECT 491.380 121.080 491.640 121.340 ;
        RECT 1076.500 121.080 1076.760 121.340 ;
      LAYER met2 ;
        RECT 493.010 500.000 493.290 504.000 ;
        RECT 493.050 498.850 493.190 500.000 ;
        RECT 492.820 498.710 493.190 498.850 ;
        RECT 492.820 488.650 492.960 498.710 ;
        RECT 492.360 488.510 492.960 488.650 ;
        RECT 492.360 472.330 492.500 488.510 ;
        RECT 491.440 472.190 492.500 472.330 ;
        RECT 491.440 121.370 491.580 472.190 ;
        RECT 491.380 121.050 491.640 121.370 ;
        RECT 1076.500 121.050 1076.760 121.370 ;
        RECT 1076.560 82.870 1076.700 121.050 ;
        RECT 1076.560 82.730 1081.760 82.870 ;
        RECT 1081.620 2.400 1081.760 82.730 ;
        RECT 1081.410 -4.800 1081.970 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 494.340 499.500 494.660 499.760 ;
        RECT 494.430 498.740 494.570 499.500 ;
        RECT 494.430 498.540 494.890 498.740 ;
        RECT 494.570 498.480 494.890 498.540 ;
      LAYER via ;
        RECT 494.370 499.500 494.630 499.760 ;
        RECT 494.600 498.480 494.860 498.740 ;
      LAYER met2 ;
        RECT 494.390 500.000 494.670 504.000 ;
        RECT 494.430 499.790 494.570 500.000 ;
        RECT 494.370 499.470 494.630 499.790 ;
        RECT 494.600 498.450 494.860 498.770 ;
        RECT 494.660 488.085 494.800 498.450 ;
        RECT 494.590 487.715 494.870 488.085 ;
        RECT 1097.190 121.875 1097.470 122.245 ;
        RECT 1097.260 17.410 1097.400 121.875 ;
        RECT 1097.260 17.270 1098.320 17.410 ;
        RECT 1098.180 2.400 1098.320 17.270 ;
        RECT 1097.970 -4.800 1098.530 2.400 ;
      LAYER via2 ;
        RECT 494.590 487.760 494.870 488.040 ;
        RECT 1097.190 121.920 1097.470 122.200 ;
      LAYER met3 ;
        RECT 494.565 488.060 494.895 488.065 ;
        RECT 494.310 488.050 494.895 488.060 ;
        RECT 494.110 487.750 494.895 488.050 ;
        RECT 494.310 487.740 494.895 487.750 ;
        RECT 494.565 487.735 494.895 487.740 ;
        RECT 494.310 122.210 494.690 122.220 ;
        RECT 1097.165 122.210 1097.495 122.225 ;
        RECT 494.310 121.910 1097.495 122.210 ;
        RECT 494.310 121.900 494.690 121.910 ;
        RECT 1097.165 121.895 1097.495 121.910 ;
      LAYER via3 ;
        RECT 494.340 487.740 494.660 488.060 ;
        RECT 494.340 121.900 494.660 122.220 ;
      LAYER met4 ;
        RECT 494.335 487.735 494.665 488.065 ;
        RECT 494.350 122.225 494.650 487.735 ;
        RECT 494.335 121.895 494.665 122.225 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 495.720 499.700 496.040 499.760 ;
        RECT 495.580 499.500 496.040 499.700 ;
        RECT 495.580 499.080 495.720 499.500 ;
        RECT 495.490 498.820 495.810 499.080 ;
      LAYER via ;
        RECT 495.750 499.500 496.010 499.760 ;
        RECT 495.520 498.820 495.780 499.080 ;
      LAYER met2 ;
        RECT 495.770 500.000 496.050 504.000 ;
        RECT 495.810 499.790 495.950 500.000 ;
        RECT 495.750 499.470 496.010 499.790 ;
        RECT 495.520 498.790 495.780 499.110 ;
        RECT 495.580 488.085 495.720 498.790 ;
        RECT 495.510 487.715 495.790 488.085 ;
        RECT 1114.670 32.795 1114.950 33.165 ;
        RECT 1114.740 2.400 1114.880 32.795 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 495.510 487.760 495.790 488.040 ;
        RECT 1114.670 32.840 1114.950 33.120 ;
      LAYER met3 ;
        RECT 495.485 488.050 495.815 488.065 ;
        RECT 496.150 488.050 496.530 488.060 ;
        RECT 495.485 487.750 496.530 488.050 ;
        RECT 495.485 487.735 495.815 487.750 ;
        RECT 496.150 487.740 496.530 487.750 ;
        RECT 496.150 33.130 496.530 33.140 ;
        RECT 1114.645 33.130 1114.975 33.145 ;
        RECT 496.150 32.830 1114.975 33.130 ;
        RECT 496.150 32.820 496.530 32.830 ;
        RECT 1114.645 32.815 1114.975 32.830 ;
      LAYER via3 ;
        RECT 496.180 487.740 496.500 488.060 ;
        RECT 496.180 32.820 496.500 33.140 ;
      LAYER met4 ;
        RECT 496.175 487.735 496.505 488.065 ;
        RECT 496.190 33.145 496.490 487.735 ;
        RECT 496.175 32.815 496.505 33.145 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.100 499.160 497.420 499.420 ;
        RECT 497.190 498.340 497.330 499.160 ;
        RECT 497.190 498.200 498.480 498.340 ;
        RECT 498.340 497.320 498.480 498.200 ;
        RECT 499.170 497.320 499.490 497.380 ;
        RECT 498.340 497.180 499.490 497.320 ;
        RECT 499.170 497.120 499.490 497.180 ;
        RECT 499.170 231.100 499.490 231.160 ;
        RECT 1125.230 231.100 1125.550 231.160 ;
        RECT 499.170 230.960 1125.550 231.100 ;
        RECT 499.170 230.900 499.490 230.960 ;
        RECT 1125.230 230.900 1125.550 230.960 ;
        RECT 1125.230 19.620 1125.550 19.680 ;
        RECT 1131.210 19.620 1131.530 19.680 ;
        RECT 1125.230 19.480 1131.530 19.620 ;
        RECT 1125.230 19.420 1125.550 19.480 ;
        RECT 1131.210 19.420 1131.530 19.480 ;
      LAYER via ;
        RECT 497.130 499.160 497.390 499.420 ;
        RECT 499.200 497.120 499.460 497.380 ;
        RECT 499.200 230.900 499.460 231.160 ;
        RECT 1125.260 230.900 1125.520 231.160 ;
        RECT 1125.260 19.420 1125.520 19.680 ;
        RECT 1131.240 19.420 1131.500 19.680 ;
      LAYER met2 ;
        RECT 497.150 500.000 497.430 504.000 ;
        RECT 497.190 499.450 497.330 500.000 ;
        RECT 497.130 499.130 497.390 499.450 ;
        RECT 499.200 497.090 499.460 497.410 ;
        RECT 499.260 231.190 499.400 497.090 ;
        RECT 499.200 230.870 499.460 231.190 ;
        RECT 1125.260 230.870 1125.520 231.190 ;
        RECT 1125.320 19.710 1125.460 230.870 ;
        RECT 1125.260 19.390 1125.520 19.710 ;
        RECT 1131.240 19.390 1131.500 19.710 ;
        RECT 1131.300 2.400 1131.440 19.390 ;
        RECT 1131.090 -4.800 1131.650 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 39.340 497.650 39.400 ;
        RECT 1147.770 39.340 1148.090 39.400 ;
        RECT 497.330 39.200 1148.090 39.340 ;
        RECT 497.330 39.140 497.650 39.200 ;
        RECT 1147.770 39.140 1148.090 39.200 ;
      LAYER via ;
        RECT 497.360 39.140 497.620 39.400 ;
        RECT 1147.800 39.140 1148.060 39.400 ;
      LAYER met2 ;
        RECT 498.530 500.000 498.810 504.000 ;
        RECT 498.570 499.645 498.710 500.000 ;
        RECT 498.500 499.275 498.780 499.645 ;
        RECT 496.430 497.915 496.710 498.285 ;
        RECT 496.500 483.070 496.640 497.915 ;
        RECT 496.500 482.930 497.100 483.070 ;
        RECT 496.960 448.570 497.100 482.930 ;
        RECT 496.960 448.430 497.560 448.570 ;
        RECT 497.420 39.430 497.560 448.430 ;
        RECT 497.360 39.110 497.620 39.430 ;
        RECT 1147.800 39.110 1148.060 39.430 ;
        RECT 1147.860 2.400 1148.000 39.110 ;
        RECT 1147.650 -4.800 1148.210 2.400 ;
      LAYER via2 ;
        RECT 498.500 499.320 498.780 499.600 ;
        RECT 496.430 497.960 496.710 498.240 ;
      LAYER met3 ;
        RECT 498.475 499.610 498.805 499.625 ;
        RECT 497.110 499.310 498.805 499.610 ;
        RECT 496.405 498.250 496.735 498.265 ;
        RECT 497.110 498.250 497.410 499.310 ;
        RECT 498.475 499.295 498.805 499.310 ;
        RECT 496.405 497.950 497.410 498.250 ;
        RECT 496.405 497.935 496.735 497.950 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.550 26.420 500.870 26.480 ;
        RECT 1164.330 26.420 1164.650 26.480 ;
        RECT 500.550 26.280 1164.650 26.420 ;
        RECT 500.550 26.220 500.870 26.280 ;
        RECT 1164.330 26.220 1164.650 26.280 ;
      LAYER via ;
        RECT 500.580 26.220 500.840 26.480 ;
        RECT 1164.360 26.220 1164.620 26.480 ;
      LAYER met2 ;
        RECT 499.910 500.000 500.190 504.000 ;
        RECT 499.950 499.645 500.090 500.000 ;
        RECT 499.880 499.275 500.160 499.645 ;
        RECT 500.570 497.915 500.850 498.285 ;
        RECT 500.640 26.510 500.780 497.915 ;
        RECT 500.580 26.190 500.840 26.510 ;
        RECT 1164.360 26.190 1164.620 26.510 ;
        RECT 1164.420 2.400 1164.560 26.190 ;
        RECT 1164.210 -4.800 1164.770 2.400 ;
      LAYER via2 ;
        RECT 499.880 499.320 500.160 499.600 ;
        RECT 500.570 497.960 500.850 498.240 ;
      LAYER met3 ;
        RECT 499.855 499.295 500.185 499.625 ;
        RECT 499.870 498.250 500.170 499.295 ;
        RECT 500.545 498.250 500.875 498.265 ;
        RECT 499.870 497.950 500.875 498.250 ;
        RECT 500.545 497.935 500.875 497.950 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 501.240 499.500 501.560 499.760 ;
        RECT 501.330 499.020 501.470 499.500 ;
        RECT 501.100 498.880 501.470 499.020 ;
        RECT 501.100 498.060 501.240 498.880 ;
        RECT 501.010 497.800 501.330 498.060 ;
      LAYER via ;
        RECT 501.270 499.500 501.530 499.760 ;
        RECT 501.040 497.800 501.300 498.060 ;
      LAYER met2 ;
        RECT 501.290 500.000 501.570 504.000 ;
        RECT 501.330 499.790 501.470 500.000 ;
        RECT 501.270 499.470 501.530 499.790 ;
        RECT 501.040 497.770 501.300 498.090 ;
        RECT 501.100 491.485 501.240 497.770 ;
        RECT 501.030 491.115 501.310 491.485 ;
        RECT 1180.910 45.715 1181.190 46.085 ;
        RECT 1180.980 2.400 1181.120 45.715 ;
        RECT 1180.770 -4.800 1181.330 2.400 ;
      LAYER via2 ;
        RECT 501.030 491.160 501.310 491.440 ;
        RECT 1180.910 45.760 1181.190 46.040 ;
      LAYER met3 ;
        RECT 499.830 491.450 500.210 491.460 ;
        RECT 501.005 491.450 501.335 491.465 ;
        RECT 499.830 491.150 501.335 491.450 ;
        RECT 499.830 491.140 500.210 491.150 ;
        RECT 501.005 491.135 501.335 491.150 ;
        RECT 499.830 46.050 500.210 46.060 ;
        RECT 1180.885 46.050 1181.215 46.065 ;
        RECT 499.830 45.750 1181.215 46.050 ;
        RECT 499.830 45.740 500.210 45.750 ;
        RECT 1180.885 45.735 1181.215 45.750 ;
      LAYER via3 ;
        RECT 499.860 491.140 500.180 491.460 ;
        RECT 499.860 45.740 500.180 46.060 ;
      LAYER met4 ;
        RECT 499.855 491.135 500.185 491.465 ;
        RECT 499.870 46.065 500.170 491.135 ;
        RECT 499.855 45.735 500.185 46.065 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.750 130.460 464.070 130.520 ;
        RECT 731.470 130.460 731.790 130.520 ;
        RECT 463.750 130.320 731.790 130.460 ;
        RECT 463.750 130.260 464.070 130.320 ;
        RECT 731.470 130.260 731.790 130.320 ;
      LAYER via ;
        RECT 463.780 130.260 464.040 130.520 ;
        RECT 731.500 130.260 731.760 130.520 ;
      LAYER met2 ;
        RECT 464.030 500.000 464.310 504.000 ;
        RECT 464.070 499.475 464.210 500.000 ;
        RECT 464.000 499.105 464.280 499.475 ;
        RECT 463.770 497.915 464.050 498.285 ;
        RECT 463.840 130.550 463.980 497.915 ;
        RECT 463.780 130.230 464.040 130.550 ;
        RECT 731.500 130.230 731.760 130.550 ;
        RECT 731.560 82.870 731.700 130.230 ;
        RECT 731.560 82.730 734.000 82.870 ;
        RECT 733.860 2.400 734.000 82.730 ;
        RECT 733.650 -4.800 734.210 2.400 ;
      LAYER via2 ;
        RECT 464.000 499.150 464.280 499.430 ;
        RECT 463.770 497.960 464.050 498.240 ;
      LAYER met3 ;
        RECT 463.975 499.125 464.305 499.455 ;
        RECT 463.990 498.265 464.290 499.125 ;
        RECT 463.745 497.950 464.290 498.265 ;
        RECT 463.745 497.935 464.075 497.950 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.670 500.000 502.950 504.000 ;
        RECT 502.710 498.680 502.850 500.000 ;
        RECT 502.710 498.540 503.080 498.680 ;
        RECT 502.940 490.805 503.080 498.540 ;
        RECT 502.870 490.435 503.150 490.805 ;
        RECT 1197.470 45.035 1197.750 45.405 ;
        RECT 1197.540 2.400 1197.680 45.035 ;
        RECT 1197.330 -4.800 1197.890 2.400 ;
      LAYER via2 ;
        RECT 502.870 490.480 503.150 490.760 ;
        RECT 1197.470 45.080 1197.750 45.360 ;
      LAYER met3 ;
        RECT 501.670 490.770 502.050 490.780 ;
        RECT 502.845 490.770 503.175 490.785 ;
        RECT 501.670 490.470 503.175 490.770 ;
        RECT 501.670 490.460 502.050 490.470 ;
        RECT 502.845 490.455 503.175 490.470 ;
        RECT 501.670 45.370 502.050 45.380 ;
        RECT 1197.445 45.370 1197.775 45.385 ;
        RECT 501.670 45.070 1197.775 45.370 ;
        RECT 501.670 45.060 502.050 45.070 ;
        RECT 1197.445 45.055 1197.775 45.070 ;
      LAYER via3 ;
        RECT 501.700 490.460 502.020 490.780 ;
        RECT 501.700 45.060 502.020 45.380 ;
      LAYER met4 ;
        RECT 501.695 490.455 502.025 490.785 ;
        RECT 501.710 45.385 502.010 490.455 ;
        RECT 501.695 45.055 502.025 45.385 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 130.120 504.550 130.180 ;
        RECT 1208.030 130.120 1208.350 130.180 ;
        RECT 504.230 129.980 1208.350 130.120 ;
        RECT 504.230 129.920 504.550 129.980 ;
        RECT 1208.030 129.920 1208.350 129.980 ;
        RECT 1208.030 19.620 1208.350 19.680 ;
        RECT 1214.010 19.620 1214.330 19.680 ;
        RECT 1208.030 19.480 1214.330 19.620 ;
        RECT 1208.030 19.420 1208.350 19.480 ;
        RECT 1214.010 19.420 1214.330 19.480 ;
      LAYER via ;
        RECT 504.260 129.920 504.520 130.180 ;
        RECT 1208.060 129.920 1208.320 130.180 ;
        RECT 1208.060 19.420 1208.320 19.680 ;
        RECT 1214.040 19.420 1214.300 19.680 ;
      LAYER met2 ;
        RECT 504.050 500.000 504.330 504.000 ;
        RECT 504.090 499.530 504.230 500.000 ;
        RECT 503.860 499.390 504.230 499.530 ;
        RECT 503.860 498.170 504.000 499.390 ;
        RECT 503.860 498.030 504.460 498.170 ;
        RECT 504.320 130.210 504.460 498.030 ;
        RECT 504.260 129.890 504.520 130.210 ;
        RECT 1208.060 129.890 1208.320 130.210 ;
        RECT 1208.120 19.710 1208.260 129.890 ;
        RECT 1208.060 19.390 1208.320 19.710 ;
        RECT 1214.040 19.390 1214.300 19.710 ;
        RECT 1214.100 2.400 1214.240 19.390 ;
        RECT 1213.890 -4.800 1214.450 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 505.380 499.500 505.700 499.760 ;
        RECT 505.470 498.400 505.610 499.500 ;
        RECT 505.470 498.200 505.930 498.400 ;
        RECT 505.610 498.140 505.930 498.200 ;
        RECT 505.610 129.780 505.930 129.840 ;
        RECT 1228.270 129.780 1228.590 129.840 ;
        RECT 505.610 129.640 1228.590 129.780 ;
        RECT 505.610 129.580 505.930 129.640 ;
        RECT 1228.270 129.580 1228.590 129.640 ;
      LAYER via ;
        RECT 505.410 499.500 505.670 499.760 ;
        RECT 505.640 498.140 505.900 498.400 ;
        RECT 505.640 129.580 505.900 129.840 ;
        RECT 1228.300 129.580 1228.560 129.840 ;
      LAYER met2 ;
        RECT 505.430 500.000 505.710 504.000 ;
        RECT 505.470 499.790 505.610 500.000 ;
        RECT 505.410 499.470 505.670 499.790 ;
        RECT 505.640 498.110 505.900 498.430 ;
        RECT 505.700 129.870 505.840 498.110 ;
        RECT 505.640 129.550 505.900 129.870 ;
        RECT 1228.300 129.550 1228.560 129.870 ;
        RECT 1228.360 82.870 1228.500 129.550 ;
        RECT 1228.360 82.730 1230.800 82.870 ;
        RECT 1230.660 2.400 1230.800 82.730 ;
        RECT 1230.450 -4.800 1231.010 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 507.910 498.340 508.230 498.400 ;
        RECT 507.080 498.200 508.230 498.340 ;
        RECT 507.080 498.060 507.220 498.200 ;
        RECT 507.910 498.140 508.230 498.200 ;
        RECT 506.990 497.800 507.310 498.060 ;
        RECT 504.690 472.840 505.010 472.900 ;
        RECT 507.910 472.840 508.230 472.900 ;
        RECT 504.690 472.700 508.230 472.840 ;
        RECT 504.690 472.640 505.010 472.700 ;
        RECT 507.910 472.640 508.230 472.700 ;
        RECT 504.690 129.440 505.010 129.500 ;
        RECT 1242.070 129.440 1242.390 129.500 ;
        RECT 504.690 129.300 1242.390 129.440 ;
        RECT 504.690 129.240 505.010 129.300 ;
        RECT 1242.070 129.240 1242.390 129.300 ;
      LAYER via ;
        RECT 507.940 498.140 508.200 498.400 ;
        RECT 507.020 497.800 507.280 498.060 ;
        RECT 504.720 472.640 504.980 472.900 ;
        RECT 507.940 472.640 508.200 472.900 ;
        RECT 504.720 129.240 504.980 129.500 ;
        RECT 1242.100 129.240 1242.360 129.500 ;
      LAYER met2 ;
        RECT 506.810 500.000 507.090 504.000 ;
        RECT 506.850 498.680 506.990 500.000 ;
        RECT 506.850 498.540 507.220 498.680 ;
        RECT 507.080 498.090 507.220 498.540 ;
        RECT 507.940 498.110 508.200 498.430 ;
        RECT 507.020 497.770 507.280 498.090 ;
        RECT 508.000 472.930 508.140 498.110 ;
        RECT 504.720 472.610 504.980 472.930 ;
        RECT 507.940 472.610 508.200 472.930 ;
        RECT 504.780 129.530 504.920 472.610 ;
        RECT 504.720 129.210 504.980 129.530 ;
        RECT 1242.100 129.210 1242.360 129.530 ;
        RECT 1242.160 82.870 1242.300 129.210 ;
        RECT 1242.160 82.730 1247.360 82.870 ;
        RECT 1247.220 2.400 1247.360 82.730 ;
        RECT 1247.010 -4.800 1247.570 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 505.150 462.640 505.470 462.700 ;
        RECT 508.370 462.640 508.690 462.700 ;
        RECT 505.150 462.500 508.690 462.640 ;
        RECT 505.150 462.440 505.470 462.500 ;
        RECT 508.370 462.440 508.690 462.500 ;
        RECT 505.150 129.100 505.470 129.160 ;
        RECT 1263.230 129.100 1263.550 129.160 ;
        RECT 505.150 128.960 1263.550 129.100 ;
        RECT 505.150 128.900 505.470 128.960 ;
        RECT 1263.230 128.900 1263.550 128.960 ;
      LAYER via ;
        RECT 505.180 462.440 505.440 462.700 ;
        RECT 508.400 462.440 508.660 462.700 ;
        RECT 505.180 128.900 505.440 129.160 ;
        RECT 1263.260 128.900 1263.520 129.160 ;
      LAYER met2 ;
        RECT 508.190 500.000 508.470 504.000 ;
        RECT 508.230 499.815 508.370 500.000 ;
        RECT 508.160 499.445 508.440 499.815 ;
        RECT 508.390 497.915 508.670 498.285 ;
        RECT 508.460 462.730 508.600 497.915 ;
        RECT 505.180 462.410 505.440 462.730 ;
        RECT 508.400 462.410 508.660 462.730 ;
        RECT 505.240 129.190 505.380 462.410 ;
        RECT 505.180 128.870 505.440 129.190 ;
        RECT 1263.260 128.870 1263.520 129.190 ;
        RECT 1263.320 82.870 1263.460 128.870 ;
        RECT 1263.320 82.730 1263.920 82.870 ;
        RECT 1263.780 2.400 1263.920 82.730 ;
        RECT 1263.570 -4.800 1264.130 2.400 ;
      LAYER via2 ;
        RECT 508.160 499.490 508.440 499.770 ;
        RECT 508.390 497.960 508.670 498.240 ;
      LAYER met3 ;
        RECT 508.135 499.610 508.465 499.795 ;
        RECT 507.230 499.465 508.465 499.610 ;
        RECT 507.230 499.310 508.450 499.465 ;
        RECT 507.230 498.250 507.530 499.310 ;
        RECT 508.365 498.250 508.695 498.265 ;
        RECT 507.230 497.950 508.695 498.250 ;
        RECT 508.365 497.935 508.695 497.950 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.570 500.000 509.850 504.000 ;
        RECT 509.610 498.680 509.750 500.000 ;
        RECT 509.610 498.540 509.980 498.680 ;
        RECT 509.840 498.285 509.980 498.540 ;
        RECT 509.770 497.915 510.050 498.285 ;
        RECT 1276.590 127.315 1276.870 127.685 ;
        RECT 1276.660 82.870 1276.800 127.315 ;
        RECT 1276.660 82.730 1280.480 82.870 ;
        RECT 1280.340 2.400 1280.480 82.730 ;
        RECT 1280.130 -4.800 1280.690 2.400 ;
      LAYER via2 ;
        RECT 509.770 497.960 510.050 498.240 ;
        RECT 1276.590 127.360 1276.870 127.640 ;
      LAYER met3 ;
        RECT 509.745 497.935 510.075 498.265 ;
        RECT 508.110 497.570 508.490 497.580 ;
        RECT 509.760 497.570 510.060 497.935 ;
        RECT 508.110 497.270 510.060 497.570 ;
        RECT 508.110 497.260 508.490 497.270 ;
        RECT 508.110 127.650 508.490 127.660 ;
        RECT 1276.565 127.650 1276.895 127.665 ;
        RECT 508.110 127.350 1276.895 127.650 ;
        RECT 508.110 127.340 508.490 127.350 ;
        RECT 1276.565 127.335 1276.895 127.350 ;
      LAYER via3 ;
        RECT 508.140 497.260 508.460 497.580 ;
        RECT 508.140 127.340 508.460 127.660 ;
      LAYER met4 ;
        RECT 508.135 497.255 508.465 497.585 ;
        RECT 508.150 127.665 508.450 497.255 ;
        RECT 508.135 127.335 508.465 127.665 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.900 499.500 511.220 499.760 ;
        RECT 510.990 496.980 511.130 499.500 ;
        RECT 514.350 496.980 514.670 497.040 ;
        RECT 510.990 496.840 514.670 496.980 ;
        RECT 514.350 496.780 514.670 496.840 ;
        RECT 514.350 135.900 514.670 135.960 ;
        RECT 1290.830 135.900 1291.150 135.960 ;
        RECT 514.350 135.760 1291.150 135.900 ;
        RECT 514.350 135.700 514.670 135.760 ;
        RECT 1290.830 135.700 1291.150 135.760 ;
        RECT 1290.830 19.620 1291.150 19.680 ;
        RECT 1296.810 19.620 1297.130 19.680 ;
        RECT 1290.830 19.480 1297.130 19.620 ;
        RECT 1290.830 19.420 1291.150 19.480 ;
        RECT 1296.810 19.420 1297.130 19.480 ;
      LAYER via ;
        RECT 510.930 499.500 511.190 499.760 ;
        RECT 514.380 496.780 514.640 497.040 ;
        RECT 514.380 135.700 514.640 135.960 ;
        RECT 1290.860 135.700 1291.120 135.960 ;
        RECT 1290.860 19.420 1291.120 19.680 ;
        RECT 1296.840 19.420 1297.100 19.680 ;
      LAYER met2 ;
        RECT 510.950 500.000 511.230 504.000 ;
        RECT 510.990 499.790 511.130 500.000 ;
        RECT 510.930 499.470 511.190 499.790 ;
        RECT 514.380 496.750 514.640 497.070 ;
        RECT 514.440 135.990 514.580 496.750 ;
        RECT 514.380 135.670 514.640 135.990 ;
        RECT 1290.860 135.670 1291.120 135.990 ;
        RECT 1290.920 19.710 1291.060 135.670 ;
        RECT 1290.860 19.390 1291.120 19.710 ;
        RECT 1296.840 19.390 1297.100 19.710 ;
        RECT 1296.900 2.400 1297.040 19.390 ;
        RECT 1296.690 -4.800 1297.250 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 512.280 499.700 512.600 499.760 ;
        RECT 512.280 499.500 512.740 499.700 ;
        RECT 512.600 497.660 512.740 499.500 ;
        RECT 513.430 497.660 513.750 497.720 ;
        RECT 512.600 497.520 513.750 497.660 ;
        RECT 513.430 497.460 513.750 497.520 ;
        RECT 513.430 135.560 513.750 135.620 ;
        RECT 1311.070 135.560 1311.390 135.620 ;
        RECT 513.430 135.420 1311.390 135.560 ;
        RECT 513.430 135.360 513.750 135.420 ;
        RECT 1311.070 135.360 1311.390 135.420 ;
      LAYER via ;
        RECT 512.310 499.500 512.570 499.760 ;
        RECT 513.460 497.460 513.720 497.720 ;
        RECT 513.460 135.360 513.720 135.620 ;
        RECT 1311.100 135.360 1311.360 135.620 ;
      LAYER met2 ;
        RECT 512.330 500.000 512.610 504.000 ;
        RECT 512.370 499.790 512.510 500.000 ;
        RECT 512.310 499.470 512.570 499.790 ;
        RECT 513.460 497.430 513.720 497.750 ;
        RECT 513.520 135.650 513.660 497.430 ;
        RECT 513.460 135.330 513.720 135.650 ;
        RECT 1311.100 135.330 1311.360 135.650 ;
        RECT 1311.160 82.870 1311.300 135.330 ;
        RECT 1311.160 82.730 1313.600 82.870 ;
        RECT 1313.460 2.400 1313.600 82.730 ;
        RECT 1313.250 -4.800 1313.810 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 513.890 135.220 514.210 135.280 ;
        RECT 1324.870 135.220 1325.190 135.280 ;
        RECT 513.890 135.080 1325.190 135.220 ;
        RECT 513.890 135.020 514.210 135.080 ;
        RECT 1324.870 135.020 1325.190 135.080 ;
      LAYER via ;
        RECT 513.920 135.020 514.180 135.280 ;
        RECT 1324.900 135.020 1325.160 135.280 ;
      LAYER met2 ;
        RECT 513.710 500.000 513.990 504.000 ;
        RECT 513.750 499.815 513.890 500.000 ;
        RECT 513.680 499.445 513.960 499.815 ;
        RECT 513.910 497.915 514.190 498.285 ;
        RECT 513.980 135.310 514.120 497.915 ;
        RECT 513.920 134.990 514.180 135.310 ;
        RECT 1324.900 134.990 1325.160 135.310 ;
        RECT 1324.960 82.870 1325.100 134.990 ;
        RECT 1324.960 82.730 1330.160 82.870 ;
        RECT 1330.020 2.400 1330.160 82.730 ;
        RECT 1329.810 -4.800 1330.370 2.400 ;
      LAYER via2 ;
        RECT 513.680 499.490 513.960 499.770 ;
        RECT 513.910 497.960 514.190 498.240 ;
      LAYER met3 ;
        RECT 513.655 499.465 513.985 499.795 ;
        RECT 513.670 498.265 513.970 499.465 ;
        RECT 513.670 497.950 514.215 498.265 ;
        RECT 513.885 497.935 514.215 497.950 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 515.040 498.820 515.360 499.080 ;
        RECT 515.130 498.400 515.270 498.820 ;
        RECT 514.810 498.200 515.270 498.400 ;
        RECT 514.810 498.140 515.130 498.200 ;
        RECT 512.050 450.740 512.370 450.800 ;
        RECT 514.810 450.740 515.130 450.800 ;
        RECT 512.050 450.600 515.130 450.740 ;
        RECT 512.050 450.540 512.370 450.600 ;
        RECT 514.810 450.540 515.130 450.600 ;
        RECT 512.050 53.620 512.370 53.680 ;
        RECT 1346.490 53.620 1346.810 53.680 ;
        RECT 512.050 53.480 1346.810 53.620 ;
        RECT 512.050 53.420 512.370 53.480 ;
        RECT 1346.490 53.420 1346.810 53.480 ;
      LAYER via ;
        RECT 515.070 498.820 515.330 499.080 ;
        RECT 514.840 498.140 515.100 498.400 ;
        RECT 512.080 450.540 512.340 450.800 ;
        RECT 514.840 450.540 515.100 450.800 ;
        RECT 512.080 53.420 512.340 53.680 ;
        RECT 1346.520 53.420 1346.780 53.680 ;
      LAYER met2 ;
        RECT 515.090 500.000 515.370 504.000 ;
        RECT 515.130 499.110 515.270 500.000 ;
        RECT 515.070 498.790 515.330 499.110 ;
        RECT 514.840 498.110 515.100 498.430 ;
        RECT 514.900 450.830 515.040 498.110 ;
        RECT 512.080 450.510 512.340 450.830 ;
        RECT 514.840 450.510 515.100 450.830 ;
        RECT 512.140 53.710 512.280 450.510 ;
        RECT 512.080 53.390 512.340 53.710 ;
        RECT 1346.520 53.390 1346.780 53.710 ;
        RECT 1346.580 2.400 1346.720 53.390 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.210 136.580 464.530 136.640 ;
        RECT 745.270 136.580 745.590 136.640 ;
        RECT 464.210 136.440 745.590 136.580 ;
        RECT 464.210 136.380 464.530 136.440 ;
        RECT 745.270 136.380 745.590 136.440 ;
      LAYER via ;
        RECT 464.240 136.380 464.500 136.640 ;
        RECT 745.300 136.380 745.560 136.640 ;
      LAYER met2 ;
        RECT 465.410 500.000 465.690 504.000 ;
        RECT 465.450 499.020 465.590 500.000 ;
        RECT 464.760 498.880 465.590 499.020 ;
        RECT 464.760 473.010 464.900 498.880 ;
        RECT 464.300 472.870 464.900 473.010 ;
        RECT 464.300 136.670 464.440 472.870 ;
        RECT 464.240 136.350 464.500 136.670 ;
        RECT 745.300 136.350 745.560 136.670 ;
        RECT 745.360 82.870 745.500 136.350 ;
        RECT 745.360 82.730 750.560 82.870 ;
        RECT 750.420 2.400 750.560 82.730 ;
        RECT 750.210 -4.800 750.770 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.420 499.500 516.740 499.760 ;
        RECT 516.510 499.080 516.650 499.500 ;
        RECT 516.420 498.820 516.740 499.080 ;
      LAYER via ;
        RECT 516.450 499.500 516.710 499.760 ;
        RECT 516.450 498.820 516.710 499.080 ;
      LAYER met2 ;
        RECT 516.470 500.000 516.750 504.000 ;
        RECT 516.510 499.790 516.650 500.000 ;
        RECT 516.450 499.470 516.710 499.790 ;
        RECT 516.450 498.965 516.710 499.110 ;
        RECT 516.440 498.595 516.720 498.965 ;
        RECT 1363.070 51.835 1363.350 52.205 ;
        RECT 1363.140 2.400 1363.280 51.835 ;
        RECT 1362.930 -4.800 1363.490 2.400 ;
      LAYER via2 ;
        RECT 516.440 498.640 516.720 498.920 ;
        RECT 1363.070 51.880 1363.350 52.160 ;
      LAYER met3 ;
        RECT 516.415 498.940 516.745 498.945 ;
        RECT 516.390 498.930 516.770 498.940 ;
        RECT 515.960 498.630 516.770 498.930 ;
        RECT 516.390 498.620 516.770 498.630 ;
        RECT 516.415 498.615 516.745 498.620 ;
        RECT 516.390 52.170 516.770 52.180 ;
        RECT 1363.045 52.170 1363.375 52.185 ;
        RECT 516.390 51.870 1363.375 52.170 ;
        RECT 516.390 51.860 516.770 51.870 ;
        RECT 1363.045 51.855 1363.375 51.870 ;
      LAYER via3 ;
        RECT 516.420 498.620 516.740 498.940 ;
        RECT 516.420 51.860 516.740 52.180 ;
      LAYER met4 ;
        RECT 516.415 498.615 516.745 498.945 ;
        RECT 516.430 52.185 516.730 498.615 ;
        RECT 516.415 51.855 516.745 52.185 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 482.700 517.890 482.760 ;
        RECT 519.410 482.700 519.730 482.760 ;
        RECT 517.570 482.560 519.730 482.700 ;
        RECT 517.570 482.500 517.890 482.560 ;
        RECT 519.410 482.500 519.730 482.560 ;
        RECT 519.410 134.880 519.730 134.940 ;
        RECT 1373.630 134.880 1373.950 134.940 ;
        RECT 519.410 134.740 1373.950 134.880 ;
        RECT 519.410 134.680 519.730 134.740 ;
        RECT 1373.630 134.680 1373.950 134.740 ;
        RECT 1373.630 19.620 1373.950 19.680 ;
        RECT 1379.610 19.620 1379.930 19.680 ;
        RECT 1373.630 19.480 1379.930 19.620 ;
        RECT 1373.630 19.420 1373.950 19.480 ;
        RECT 1379.610 19.420 1379.930 19.480 ;
      LAYER via ;
        RECT 517.600 482.500 517.860 482.760 ;
        RECT 519.440 482.500 519.700 482.760 ;
        RECT 519.440 134.680 519.700 134.940 ;
        RECT 1373.660 134.680 1373.920 134.940 ;
        RECT 1373.660 19.420 1373.920 19.680 ;
        RECT 1379.640 19.420 1379.900 19.680 ;
      LAYER met2 ;
        RECT 517.850 500.000 518.130 504.000 ;
        RECT 517.890 499.645 518.030 500.000 ;
        RECT 517.820 499.275 518.100 499.645 ;
        RECT 517.590 497.915 517.870 498.285 ;
        RECT 517.660 482.790 517.800 497.915 ;
        RECT 517.600 482.470 517.860 482.790 ;
        RECT 519.440 482.470 519.700 482.790 ;
        RECT 519.500 134.970 519.640 482.470 ;
        RECT 519.440 134.650 519.700 134.970 ;
        RECT 1373.660 134.650 1373.920 134.970 ;
        RECT 1373.720 19.710 1373.860 134.650 ;
        RECT 1373.660 19.390 1373.920 19.710 ;
        RECT 1379.640 19.390 1379.900 19.710 ;
        RECT 1379.700 2.400 1379.840 19.390 ;
        RECT 1379.490 -4.800 1380.050 2.400 ;
      LAYER via2 ;
        RECT 517.820 499.320 518.100 499.600 ;
        RECT 517.590 497.960 517.870 498.240 ;
      LAYER met3 ;
        RECT 517.795 499.610 518.125 499.625 ;
        RECT 517.120 499.310 518.125 499.610 ;
        RECT 517.120 498.930 517.420 499.310 ;
        RECT 517.795 499.295 518.125 499.310 ;
        RECT 517.120 498.630 517.650 498.930 ;
        RECT 517.350 498.265 517.650 498.630 ;
        RECT 517.350 497.950 517.895 498.265 ;
        RECT 517.565 497.935 517.895 497.950 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.180 499.500 519.500 499.760 ;
        RECT 519.270 498.740 519.410 499.500 ;
        RECT 519.270 498.540 519.730 498.740 ;
        RECT 519.410 498.480 519.730 498.540 ;
        RECT 518.950 134.540 519.270 134.600 ;
        RECT 1393.870 134.540 1394.190 134.600 ;
        RECT 518.950 134.400 1394.190 134.540 ;
        RECT 518.950 134.340 519.270 134.400 ;
        RECT 1393.870 134.340 1394.190 134.400 ;
      LAYER via ;
        RECT 519.210 499.500 519.470 499.760 ;
        RECT 519.440 498.480 519.700 498.740 ;
        RECT 518.980 134.340 519.240 134.600 ;
        RECT 1393.900 134.340 1394.160 134.600 ;
      LAYER met2 ;
        RECT 519.230 500.000 519.510 504.000 ;
        RECT 519.270 499.790 519.410 500.000 ;
        RECT 519.210 499.470 519.470 499.790 ;
        RECT 519.440 498.450 519.700 498.770 ;
        RECT 519.500 483.070 519.640 498.450 ;
        RECT 519.040 482.930 519.640 483.070 ;
        RECT 519.040 134.630 519.180 482.930 ;
        RECT 518.980 134.310 519.240 134.630 ;
        RECT 1393.900 134.310 1394.160 134.630 ;
        RECT 1393.960 82.870 1394.100 134.310 ;
        RECT 1393.960 82.730 1396.400 82.870 ;
        RECT 1396.260 2.400 1396.400 82.730 ;
        RECT 1396.050 -4.800 1396.610 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.560 499.500 520.880 499.760 ;
        RECT 520.650 498.400 520.790 499.500 ;
        RECT 520.330 498.200 520.790 498.400 ;
        RECT 520.330 498.140 520.650 498.200 ;
        RECT 520.790 142.700 521.110 142.760 ;
        RECT 1407.670 142.700 1407.990 142.760 ;
        RECT 520.790 142.560 1407.990 142.700 ;
        RECT 520.790 142.500 521.110 142.560 ;
        RECT 1407.670 142.500 1407.990 142.560 ;
      LAYER via ;
        RECT 520.590 499.500 520.850 499.760 ;
        RECT 520.360 498.140 520.620 498.400 ;
        RECT 520.820 142.500 521.080 142.760 ;
        RECT 1407.700 142.500 1407.960 142.760 ;
      LAYER met2 ;
        RECT 520.610 500.000 520.890 504.000 ;
        RECT 520.650 499.790 520.790 500.000 ;
        RECT 520.590 499.470 520.850 499.790 ;
        RECT 520.360 498.110 520.620 498.430 ;
        RECT 520.420 478.280 520.560 498.110 ;
        RECT 520.420 478.140 521.020 478.280 ;
        RECT 520.880 142.790 521.020 478.140 ;
        RECT 520.820 142.470 521.080 142.790 ;
        RECT 1407.700 142.470 1407.960 142.790 ;
        RECT 1407.760 82.870 1407.900 142.470 ;
        RECT 1407.760 82.730 1412.960 82.870 ;
        RECT 1412.820 2.400 1412.960 82.730 ;
        RECT 1412.610 -4.800 1413.170 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.940 499.500 522.260 499.760 ;
        RECT 522.030 498.400 522.170 499.500 ;
        RECT 522.030 498.200 522.490 498.400 ;
        RECT 522.170 498.140 522.490 498.200 ;
      LAYER via ;
        RECT 521.970 499.500 522.230 499.760 ;
        RECT 522.200 498.140 522.460 498.400 ;
      LAYER met2 ;
        RECT 521.990 500.000 522.270 504.000 ;
        RECT 522.030 499.790 522.170 500.000 ;
        RECT 521.970 499.470 522.230 499.790 ;
        RECT 522.200 498.110 522.460 498.430 ;
        RECT 522.260 478.565 522.400 498.110 ;
        RECT 522.190 478.195 522.470 478.565 ;
        RECT 1428.850 141.595 1429.130 141.965 ;
        RECT 1428.920 82.870 1429.060 141.595 ;
        RECT 1428.920 82.730 1429.520 82.870 ;
        RECT 1429.380 2.400 1429.520 82.730 ;
        RECT 1429.170 -4.800 1429.730 2.400 ;
      LAYER via2 ;
        RECT 522.190 478.240 522.470 478.520 ;
        RECT 1428.850 141.640 1429.130 141.920 ;
      LAYER met3 ;
        RECT 522.165 478.530 522.495 478.545 ;
        RECT 522.830 478.530 523.210 478.540 ;
        RECT 522.165 478.230 523.210 478.530 ;
        RECT 522.165 478.215 522.495 478.230 ;
        RECT 522.830 478.220 523.210 478.230 ;
        RECT 522.830 141.930 523.210 141.940 ;
        RECT 1428.825 141.930 1429.155 141.945 ;
        RECT 522.830 141.630 1429.155 141.930 ;
        RECT 522.830 141.620 523.210 141.630 ;
        RECT 1428.825 141.615 1429.155 141.630 ;
      LAYER via3 ;
        RECT 522.860 478.220 523.180 478.540 ;
        RECT 522.860 141.620 523.180 141.940 ;
      LAYER met4 ;
        RECT 522.855 478.215 523.185 478.545 ;
        RECT 522.870 141.945 523.170 478.215 ;
        RECT 522.855 141.615 523.185 141.945 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.570 499.900 523.550 500.040 ;
        RECT 521.570 497.040 521.710 499.900 ;
        RECT 523.410 499.760 523.550 499.900 ;
        RECT 523.320 499.500 523.640 499.760 ;
        RECT 521.250 496.840 521.710 497.040 ;
        RECT 521.250 496.780 521.570 496.840 ;
      LAYER via ;
        RECT 523.350 499.500 523.610 499.760 ;
        RECT 521.280 496.780 521.540 497.040 ;
      LAYER met2 ;
        RECT 523.370 500.000 523.650 504.000 ;
        RECT 523.410 499.790 523.550 500.000 ;
        RECT 523.350 499.470 523.610 499.790 ;
        RECT 521.280 496.750 521.540 497.070 ;
        RECT 521.340 482.645 521.480 496.750 ;
        RECT 521.270 482.275 521.550 482.645 ;
        RECT 1445.870 51.155 1446.150 51.525 ;
        RECT 1445.940 2.400 1446.080 51.155 ;
        RECT 1445.730 -4.800 1446.290 2.400 ;
      LAYER via2 ;
        RECT 521.270 482.320 521.550 482.600 ;
        RECT 1445.870 51.200 1446.150 51.480 ;
      LAYER met3 ;
        RECT 521.245 482.620 521.575 482.625 ;
        RECT 520.990 482.610 521.575 482.620 ;
        RECT 520.790 482.310 521.575 482.610 ;
        RECT 520.990 482.300 521.575 482.310 ;
        RECT 521.245 482.295 521.575 482.300 ;
        RECT 520.990 51.490 521.370 51.500 ;
        RECT 1445.845 51.490 1446.175 51.505 ;
        RECT 520.990 51.190 1446.175 51.490 ;
        RECT 520.990 51.180 521.370 51.190 ;
        RECT 1445.845 51.175 1446.175 51.190 ;
      LAYER via3 ;
        RECT 521.020 482.300 521.340 482.620 ;
        RECT 521.020 51.180 521.340 51.500 ;
      LAYER met4 ;
        RECT 521.015 482.295 521.345 482.625 ;
        RECT 521.030 51.505 521.330 482.295 ;
        RECT 521.015 51.175 521.345 51.505 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 478.620 525.250 478.680 ;
        RECT 526.770 478.620 527.090 478.680 ;
        RECT 524.930 478.480 527.090 478.620 ;
        RECT 524.930 478.420 525.250 478.480 ;
        RECT 526.770 478.420 527.090 478.480 ;
        RECT 526.770 142.360 527.090 142.420 ;
        RECT 1456.430 142.360 1456.750 142.420 ;
        RECT 526.770 142.220 1456.750 142.360 ;
        RECT 526.770 142.160 527.090 142.220 ;
        RECT 1456.430 142.160 1456.750 142.220 ;
        RECT 1456.430 19.960 1456.750 20.020 ;
        RECT 1462.410 19.960 1462.730 20.020 ;
        RECT 1456.430 19.820 1462.730 19.960 ;
        RECT 1456.430 19.760 1456.750 19.820 ;
        RECT 1462.410 19.760 1462.730 19.820 ;
      LAYER via ;
        RECT 524.960 478.420 525.220 478.680 ;
        RECT 526.800 478.420 527.060 478.680 ;
        RECT 526.800 142.160 527.060 142.420 ;
        RECT 1456.460 142.160 1456.720 142.420 ;
        RECT 1456.460 19.760 1456.720 20.020 ;
        RECT 1462.440 19.760 1462.700 20.020 ;
      LAYER met2 ;
        RECT 524.750 500.000 525.030 504.000 ;
        RECT 524.790 499.815 524.930 500.000 ;
        RECT 524.720 499.445 525.000 499.815 ;
        RECT 524.950 498.595 525.230 498.965 ;
        RECT 525.020 478.710 525.160 498.595 ;
        RECT 524.960 478.390 525.220 478.710 ;
        RECT 526.800 478.390 527.060 478.710 ;
        RECT 526.860 142.450 527.000 478.390 ;
        RECT 526.800 142.130 527.060 142.450 ;
        RECT 1456.460 142.130 1456.720 142.450 ;
        RECT 1456.520 20.050 1456.660 142.130 ;
        RECT 1456.460 19.730 1456.720 20.050 ;
        RECT 1462.440 19.730 1462.700 20.050 ;
        RECT 1462.500 2.400 1462.640 19.730 ;
        RECT 1462.290 -4.800 1462.850 2.400 ;
      LAYER via2 ;
        RECT 524.720 499.490 525.000 499.770 ;
        RECT 524.950 498.640 525.230 498.920 ;
      LAYER met3 ;
        RECT 524.695 499.465 525.025 499.795 ;
        RECT 524.710 498.945 525.010 499.465 ;
        RECT 524.710 498.630 525.255 498.945 ;
        RECT 524.925 498.615 525.255 498.630 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.850 485.080 526.170 485.140 ;
        RECT 527.230 485.080 527.550 485.140 ;
        RECT 525.850 484.940 527.550 485.080 ;
        RECT 525.850 484.880 526.170 484.940 ;
        RECT 527.230 484.880 527.550 484.940 ;
        RECT 527.230 142.020 527.550 142.080 ;
        RECT 1476.670 142.020 1476.990 142.080 ;
        RECT 527.230 141.880 1476.990 142.020 ;
        RECT 527.230 141.820 527.550 141.880 ;
        RECT 1476.670 141.820 1476.990 141.880 ;
      LAYER via ;
        RECT 525.880 484.880 526.140 485.140 ;
        RECT 527.260 484.880 527.520 485.140 ;
        RECT 527.260 141.820 527.520 142.080 ;
        RECT 1476.700 141.820 1476.960 142.080 ;
      LAYER met2 ;
        RECT 526.130 500.000 526.410 504.000 ;
        RECT 526.170 497.660 526.310 500.000 ;
        RECT 525.940 497.520 526.310 497.660 ;
        RECT 525.940 485.170 526.080 497.520 ;
        RECT 525.880 484.850 526.140 485.170 ;
        RECT 527.260 484.850 527.520 485.170 ;
        RECT 527.320 142.110 527.460 484.850 ;
        RECT 527.260 141.790 527.520 142.110 ;
        RECT 1476.700 141.790 1476.960 142.110 ;
        RECT 1476.760 82.870 1476.900 141.790 ;
        RECT 1476.760 82.730 1479.200 82.870 ;
        RECT 1479.060 2.400 1479.200 82.730 ;
        RECT 1478.850 -4.800 1479.410 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.460 499.500 527.780 499.760 ;
        RECT 527.550 498.400 527.690 499.500 ;
        RECT 527.550 498.200 528.010 498.400 ;
        RECT 527.690 498.140 528.010 498.200 ;
        RECT 524.470 486.440 524.790 486.500 ;
        RECT 527.690 486.440 528.010 486.500 ;
        RECT 524.470 486.300 528.010 486.440 ;
        RECT 524.470 486.240 524.790 486.300 ;
        RECT 527.690 486.240 528.010 486.300 ;
        RECT 524.470 26.080 524.790 26.140 ;
        RECT 1495.530 26.080 1495.850 26.140 ;
        RECT 524.470 25.940 1495.850 26.080 ;
        RECT 524.470 25.880 524.790 25.940 ;
        RECT 1495.530 25.880 1495.850 25.940 ;
      LAYER via ;
        RECT 527.490 499.500 527.750 499.760 ;
        RECT 527.720 498.140 527.980 498.400 ;
        RECT 524.500 486.240 524.760 486.500 ;
        RECT 527.720 486.240 527.980 486.500 ;
        RECT 524.500 25.880 524.760 26.140 ;
        RECT 1495.560 25.880 1495.820 26.140 ;
      LAYER met2 ;
        RECT 527.510 500.000 527.790 504.000 ;
        RECT 527.550 499.790 527.690 500.000 ;
        RECT 527.490 499.470 527.750 499.790 ;
        RECT 527.720 498.110 527.980 498.430 ;
        RECT 527.780 486.530 527.920 498.110 ;
        RECT 524.500 486.210 524.760 486.530 ;
        RECT 527.720 486.210 527.980 486.530 ;
        RECT 524.560 26.170 524.700 486.210 ;
        RECT 524.500 25.850 524.760 26.170 ;
        RECT 1495.560 25.850 1495.820 26.170 ;
        RECT 1495.620 2.400 1495.760 25.850 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.690 204.920 528.010 204.980 ;
        RECT 1511.630 204.920 1511.950 204.980 ;
        RECT 527.690 204.780 1511.950 204.920 ;
        RECT 527.690 204.720 528.010 204.780 ;
        RECT 1511.630 204.720 1511.950 204.780 ;
      LAYER via ;
        RECT 527.720 204.720 527.980 204.980 ;
        RECT 1511.660 204.720 1511.920 204.980 ;
      LAYER met2 ;
        RECT 528.890 500.000 529.170 504.000 ;
        RECT 528.930 498.340 529.070 500.000 ;
        RECT 528.700 498.200 529.070 498.340 ;
        RECT 528.700 483.890 528.840 498.200 ;
        RECT 527.780 483.750 528.840 483.890 ;
        RECT 527.780 205.010 527.920 483.750 ;
        RECT 527.720 204.690 527.980 205.010 ;
        RECT 1511.660 204.690 1511.920 205.010 ;
        RECT 1511.720 82.870 1511.860 204.690 ;
        RECT 1511.720 82.730 1512.320 82.870 ;
        RECT 1512.180 2.400 1512.320 82.730 ;
        RECT 1511.970 -4.800 1512.530 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.740 499.500 467.060 499.760 ;
        RECT 466.830 499.080 466.970 499.500 ;
        RECT 466.510 498.880 466.970 499.080 ;
        RECT 466.510 498.820 466.830 498.880 ;
      LAYER via ;
        RECT 466.770 499.500 467.030 499.760 ;
        RECT 466.540 498.820 466.800 499.080 ;
      LAYER met2 ;
        RECT 466.790 500.000 467.070 504.000 ;
        RECT 466.830 499.790 466.970 500.000 ;
        RECT 466.770 499.470 467.030 499.790 ;
        RECT 466.540 498.790 466.800 499.110 ;
        RECT 466.600 498.285 466.740 498.790 ;
        RECT 466.530 497.915 466.810 498.285 ;
        RECT 766.450 142.275 766.730 142.645 ;
        RECT 766.520 82.870 766.660 142.275 ;
        RECT 766.520 82.730 767.120 82.870 ;
        RECT 766.980 2.400 767.120 82.730 ;
        RECT 766.770 -4.800 767.330 2.400 ;
      LAYER via2 ;
        RECT 466.530 497.960 466.810 498.240 ;
        RECT 766.450 142.320 766.730 142.600 ;
      LAYER met3 ;
        RECT 466.505 498.250 466.835 498.265 ;
        RECT 467.630 498.250 468.010 498.260 ;
        RECT 466.505 497.950 468.010 498.250 ;
        RECT 466.505 497.935 466.835 497.950 ;
        RECT 467.630 497.940 468.010 497.950 ;
        RECT 467.630 142.610 468.010 142.620 ;
        RECT 766.425 142.610 766.755 142.625 ;
        RECT 467.630 142.310 766.755 142.610 ;
        RECT 467.630 142.300 468.010 142.310 ;
        RECT 766.425 142.295 766.755 142.310 ;
      LAYER via3 ;
        RECT 467.660 497.940 467.980 498.260 ;
        RECT 467.660 142.300 467.980 142.620 ;
      LAYER met4 ;
        RECT 467.655 497.935 467.985 498.265 ;
        RECT 467.670 142.625 467.970 497.935 ;
        RECT 467.655 142.295 467.985 142.625 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.270 500.000 530.550 504.000 ;
        RECT 530.310 499.815 530.450 500.000 ;
        RECT 530.240 499.445 530.520 499.815 ;
        RECT 1524.990 423.795 1525.270 424.165 ;
        RECT 1525.060 82.870 1525.200 423.795 ;
        RECT 1525.060 82.730 1528.880 82.870 ;
        RECT 1528.740 2.400 1528.880 82.730 ;
        RECT 1528.530 -4.800 1529.090 2.400 ;
      LAYER via2 ;
        RECT 530.240 499.490 530.520 499.770 ;
        RECT 1524.990 423.840 1525.270 424.120 ;
      LAYER met3 ;
        RECT 530.215 499.620 530.545 499.795 ;
        RECT 530.190 499.610 530.570 499.620 ;
        RECT 530.190 499.310 530.830 499.610 ;
        RECT 530.190 499.300 530.570 499.310 ;
        RECT 530.190 424.130 530.570 424.140 ;
        RECT 1524.965 424.130 1525.295 424.145 ;
        RECT 530.190 423.830 1525.295 424.130 ;
        RECT 530.190 423.820 530.570 423.830 ;
        RECT 1524.965 423.815 1525.295 423.830 ;
      LAYER via3 ;
        RECT 530.220 499.300 530.540 499.620 ;
        RECT 530.220 423.820 530.540 424.140 ;
      LAYER met4 ;
        RECT 530.215 499.295 530.545 499.625 ;
        RECT 530.230 424.145 530.530 499.295 ;
        RECT 530.215 423.815 530.545 424.145 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.600 499.500 531.920 499.760 ;
        RECT 531.690 498.740 531.830 499.500 ;
        RECT 531.370 498.540 531.830 498.740 ;
        RECT 531.370 498.480 531.690 498.540 ;
        RECT 531.370 483.040 531.690 483.100 ;
        RECT 533.670 483.040 533.990 483.100 ;
        RECT 531.370 482.900 533.990 483.040 ;
        RECT 531.370 482.840 531.690 482.900 ;
        RECT 533.670 482.840 533.990 482.900 ;
        RECT 533.670 150.520 533.990 150.580 ;
        RECT 1539.230 150.520 1539.550 150.580 ;
        RECT 533.670 150.380 1539.550 150.520 ;
        RECT 533.670 150.320 533.990 150.380 ;
        RECT 1539.230 150.320 1539.550 150.380 ;
        RECT 1539.230 20.300 1539.550 20.360 ;
        RECT 1545.210 20.300 1545.530 20.360 ;
        RECT 1539.230 20.160 1545.530 20.300 ;
        RECT 1539.230 20.100 1539.550 20.160 ;
        RECT 1545.210 20.100 1545.530 20.160 ;
      LAYER via ;
        RECT 531.630 499.500 531.890 499.760 ;
        RECT 531.400 498.480 531.660 498.740 ;
        RECT 531.400 482.840 531.660 483.100 ;
        RECT 533.700 482.840 533.960 483.100 ;
        RECT 533.700 150.320 533.960 150.580 ;
        RECT 1539.260 150.320 1539.520 150.580 ;
        RECT 1539.260 20.100 1539.520 20.360 ;
        RECT 1545.240 20.100 1545.500 20.360 ;
      LAYER met2 ;
        RECT 531.650 500.000 531.930 504.000 ;
        RECT 531.690 499.790 531.830 500.000 ;
        RECT 531.630 499.470 531.890 499.790 ;
        RECT 531.400 498.450 531.660 498.770 ;
        RECT 531.460 483.130 531.600 498.450 ;
        RECT 531.400 482.810 531.660 483.130 ;
        RECT 533.700 482.810 533.960 483.130 ;
        RECT 533.760 150.610 533.900 482.810 ;
        RECT 533.700 150.290 533.960 150.610 ;
        RECT 1539.260 150.290 1539.520 150.610 ;
        RECT 1539.320 20.390 1539.460 150.290 ;
        RECT 1539.260 20.070 1539.520 20.390 ;
        RECT 1545.240 20.070 1545.500 20.390 ;
        RECT 1545.300 2.400 1545.440 20.070 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.750 149.840 533.070 149.900 ;
        RECT 1559.470 149.840 1559.790 149.900 ;
        RECT 532.750 149.700 1559.790 149.840 ;
        RECT 532.750 149.640 533.070 149.700 ;
        RECT 1559.470 149.640 1559.790 149.700 ;
      LAYER via ;
        RECT 532.780 149.640 533.040 149.900 ;
        RECT 1559.500 149.640 1559.760 149.900 ;
      LAYER met2 ;
        RECT 533.030 500.000 533.310 504.000 ;
        RECT 533.070 498.680 533.210 500.000 ;
        RECT 532.840 498.540 533.210 498.680 ;
        RECT 532.840 149.930 532.980 498.540 ;
        RECT 532.780 149.610 533.040 149.930 ;
        RECT 1559.500 149.610 1559.760 149.930 ;
        RECT 1559.560 82.870 1559.700 149.610 ;
        RECT 1559.560 82.730 1562.000 82.870 ;
        RECT 1561.860 2.400 1562.000 82.730 ;
        RECT 1561.650 -4.800 1562.210 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.360 499.700 534.680 499.760 ;
        RECT 533.990 499.560 534.680 499.700 ;
        RECT 533.990 497.720 534.130 499.560 ;
        RECT 534.360 499.500 534.680 499.560 ;
        RECT 533.670 497.520 534.130 497.720 ;
        RECT 533.670 497.460 533.990 497.520 ;
        RECT 532.290 149.160 532.610 149.220 ;
        RECT 1573.270 149.160 1573.590 149.220 ;
        RECT 532.290 149.020 1573.590 149.160 ;
        RECT 532.290 148.960 532.610 149.020 ;
        RECT 1573.270 148.960 1573.590 149.020 ;
      LAYER via ;
        RECT 534.390 499.500 534.650 499.760 ;
        RECT 533.700 497.460 533.960 497.720 ;
        RECT 532.320 148.960 532.580 149.220 ;
        RECT 1573.300 148.960 1573.560 149.220 ;
      LAYER met2 ;
        RECT 534.410 500.000 534.690 504.000 ;
        RECT 534.450 499.790 534.590 500.000 ;
        RECT 534.390 499.470 534.650 499.790 ;
        RECT 533.700 497.430 533.960 497.750 ;
        RECT 533.760 484.005 533.900 497.430 ;
        RECT 533.690 483.635 533.970 484.005 ;
        RECT 532.310 482.955 532.590 483.325 ;
        RECT 532.380 149.250 532.520 482.955 ;
        RECT 532.320 148.930 532.580 149.250 ;
        RECT 1573.300 148.930 1573.560 149.250 ;
        RECT 1573.360 82.870 1573.500 148.930 ;
        RECT 1573.360 82.730 1578.560 82.870 ;
        RECT 1578.420 2.400 1578.560 82.730 ;
        RECT 1578.210 -4.800 1578.770 2.400 ;
      LAYER via2 ;
        RECT 533.690 483.680 533.970 483.960 ;
        RECT 532.310 483.000 532.590 483.280 ;
      LAYER met3 ;
        RECT 533.665 483.970 533.995 483.985 ;
        RECT 532.300 483.670 533.995 483.970 ;
        RECT 532.300 483.305 532.600 483.670 ;
        RECT 533.665 483.655 533.995 483.670 ;
        RECT 532.285 482.975 532.615 483.305 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 479.300 531.690 479.360 ;
        RECT 535.970 479.300 536.290 479.360 ;
        RECT 531.370 479.160 536.290 479.300 ;
        RECT 531.370 479.100 531.690 479.160 ;
        RECT 535.970 479.100 536.290 479.160 ;
        RECT 531.370 60.420 531.690 60.480 ;
        RECT 1594.890 60.420 1595.210 60.480 ;
        RECT 531.370 60.280 1595.210 60.420 ;
        RECT 531.370 60.220 531.690 60.280 ;
        RECT 1594.890 60.220 1595.210 60.280 ;
      LAYER via ;
        RECT 531.400 479.100 531.660 479.360 ;
        RECT 536.000 479.100 536.260 479.360 ;
        RECT 531.400 60.220 531.660 60.480 ;
        RECT 1594.920 60.220 1595.180 60.480 ;
      LAYER met2 ;
        RECT 535.790 500.000 536.070 504.000 ;
        RECT 535.830 498.680 535.970 500.000 ;
        RECT 535.600 498.540 535.970 498.680 ;
        RECT 535.600 496.870 535.740 498.540 ;
        RECT 535.600 496.730 536.200 496.870 ;
        RECT 536.060 479.390 536.200 496.730 ;
        RECT 531.400 479.070 531.660 479.390 ;
        RECT 536.000 479.070 536.260 479.390 ;
        RECT 531.460 60.510 531.600 479.070 ;
        RECT 531.400 60.190 531.660 60.510 ;
        RECT 1594.920 60.190 1595.180 60.510 ;
        RECT 1594.980 2.400 1595.120 60.190 ;
        RECT 1594.770 -4.800 1595.330 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.170 500.000 537.450 504.000 ;
        RECT 537.210 499.700 537.350 500.000 ;
        RECT 536.980 499.645 537.350 499.700 ;
        RECT 536.910 499.560 537.350 499.645 ;
        RECT 536.910 499.275 537.190 499.560 ;
        RECT 1611.470 66.115 1611.750 66.485 ;
        RECT 1611.540 2.400 1611.680 66.115 ;
        RECT 1611.330 -4.800 1611.890 2.400 ;
      LAYER via2 ;
        RECT 536.910 499.320 537.190 499.600 ;
        RECT 1611.470 66.160 1611.750 66.440 ;
      LAYER met3 ;
        RECT 536.885 499.620 537.215 499.625 ;
        RECT 536.630 499.610 537.215 499.620 ;
        RECT 536.430 499.310 537.215 499.610 ;
        RECT 536.630 499.300 537.215 499.310 ;
        RECT 536.885 499.295 537.215 499.300 ;
        RECT 536.630 66.450 537.010 66.460 ;
        RECT 1611.445 66.450 1611.775 66.465 ;
        RECT 536.630 66.150 1611.775 66.450 ;
        RECT 536.630 66.140 537.010 66.150 ;
        RECT 1611.445 66.135 1611.775 66.150 ;
      LAYER via3 ;
        RECT 536.660 499.300 536.980 499.620 ;
        RECT 536.660 66.140 536.980 66.460 ;
      LAYER met4 ;
        RECT 536.655 499.295 536.985 499.625 ;
        RECT 536.670 66.465 536.970 499.295 ;
        RECT 536.655 66.135 536.985 66.465 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.500 499.700 538.820 499.760 ;
        RECT 538.500 499.500 538.960 499.700 ;
        RECT 536.890 498.000 537.210 498.060 ;
        RECT 538.820 498.000 538.960 499.500 ;
        RECT 536.890 497.860 538.960 498.000 ;
        RECT 536.890 497.800 537.210 497.860 ;
        RECT 536.890 480.660 537.210 480.720 ;
        RECT 539.650 480.660 539.970 480.720 ;
        RECT 536.890 480.520 539.970 480.660 ;
        RECT 536.890 480.460 537.210 480.520 ;
        RECT 539.650 480.460 539.970 480.520 ;
        RECT 540.570 148.820 540.890 148.880 ;
        RECT 1622.030 148.820 1622.350 148.880 ;
        RECT 540.570 148.680 1622.350 148.820 ;
        RECT 540.570 148.620 540.890 148.680 ;
        RECT 1622.030 148.620 1622.350 148.680 ;
        RECT 1622.030 20.300 1622.350 20.360 ;
        RECT 1628.010 20.300 1628.330 20.360 ;
        RECT 1622.030 20.160 1628.330 20.300 ;
        RECT 1622.030 20.100 1622.350 20.160 ;
        RECT 1628.010 20.100 1628.330 20.160 ;
      LAYER via ;
        RECT 538.530 499.500 538.790 499.760 ;
        RECT 536.920 497.800 537.180 498.060 ;
        RECT 536.920 480.460 537.180 480.720 ;
        RECT 539.680 480.460 539.940 480.720 ;
        RECT 540.600 148.620 540.860 148.880 ;
        RECT 1622.060 148.620 1622.320 148.880 ;
        RECT 1622.060 20.100 1622.320 20.360 ;
        RECT 1628.040 20.100 1628.300 20.360 ;
      LAYER met2 ;
        RECT 538.550 500.000 538.830 504.000 ;
        RECT 538.590 499.790 538.730 500.000 ;
        RECT 538.530 499.470 538.790 499.790 ;
        RECT 536.920 497.770 537.180 498.090 ;
        RECT 536.980 480.750 537.120 497.770 ;
        RECT 536.920 480.430 537.180 480.750 ;
        RECT 539.680 480.430 539.940 480.750 ;
        RECT 539.740 451.930 539.880 480.430 ;
        RECT 539.740 451.790 540.800 451.930 ;
        RECT 540.660 148.910 540.800 451.790 ;
        RECT 540.600 148.590 540.860 148.910 ;
        RECT 1622.060 148.590 1622.320 148.910 ;
        RECT 1622.120 20.390 1622.260 148.590 ;
        RECT 1622.060 20.070 1622.320 20.390 ;
        RECT 1628.040 20.070 1628.300 20.390 ;
        RECT 1628.100 2.400 1628.240 20.070 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.880 499.500 540.200 499.760 ;
        RECT 539.970 498.000 540.110 499.500 ;
        RECT 540.570 498.000 540.890 498.060 ;
        RECT 539.970 497.860 540.890 498.000 ;
        RECT 540.570 497.800 540.890 497.860 ;
        RECT 541.030 148.480 541.350 148.540 ;
        RECT 1642.270 148.480 1642.590 148.540 ;
        RECT 541.030 148.340 1642.590 148.480 ;
        RECT 541.030 148.280 541.350 148.340 ;
        RECT 1642.270 148.280 1642.590 148.340 ;
      LAYER via ;
        RECT 539.910 499.500 540.170 499.760 ;
        RECT 540.600 497.800 540.860 498.060 ;
        RECT 541.060 148.280 541.320 148.540 ;
        RECT 1642.300 148.280 1642.560 148.540 ;
      LAYER met2 ;
        RECT 539.930 500.000 540.210 504.000 ;
        RECT 539.970 499.790 540.110 500.000 ;
        RECT 539.910 499.470 540.170 499.790 ;
        RECT 540.600 497.770 540.860 498.090 ;
        RECT 540.660 455.470 540.800 497.770 ;
        RECT 540.660 455.330 541.260 455.470 ;
        RECT 541.120 148.570 541.260 455.330 ;
        RECT 541.060 148.250 541.320 148.570 ;
        RECT 1642.300 148.250 1642.560 148.570 ;
        RECT 1642.360 82.870 1642.500 148.250 ;
        RECT 1642.360 82.730 1644.800 82.870 ;
        RECT 1644.660 2.400 1644.800 82.730 ;
        RECT 1644.450 -4.800 1645.010 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.650 451.420 539.970 451.480 ;
        RECT 541.490 451.420 541.810 451.480 ;
        RECT 539.650 451.280 541.810 451.420 ;
        RECT 539.650 451.220 539.970 451.280 ;
        RECT 541.490 451.220 541.810 451.280 ;
        RECT 539.650 67.220 539.970 67.280 ;
        RECT 1661.130 67.220 1661.450 67.280 ;
        RECT 539.650 67.080 1661.450 67.220 ;
        RECT 539.650 67.020 539.970 67.080 ;
        RECT 1661.130 67.020 1661.450 67.080 ;
      LAYER via ;
        RECT 539.680 451.220 539.940 451.480 ;
        RECT 541.520 451.220 541.780 451.480 ;
        RECT 539.680 67.020 539.940 67.280 ;
        RECT 1661.160 67.020 1661.420 67.280 ;
      LAYER met2 ;
        RECT 541.310 500.000 541.590 504.000 ;
        RECT 541.350 499.815 541.490 500.000 ;
        RECT 541.280 499.445 541.560 499.815 ;
        RECT 541.510 497.915 541.790 498.285 ;
        RECT 541.580 451.510 541.720 497.915 ;
        RECT 539.680 451.190 539.940 451.510 ;
        RECT 541.520 451.190 541.780 451.510 ;
        RECT 539.740 67.310 539.880 451.190 ;
        RECT 539.680 66.990 539.940 67.310 ;
        RECT 1661.160 66.990 1661.420 67.310 ;
        RECT 1661.220 2.400 1661.360 66.990 ;
        RECT 1661.010 -4.800 1661.570 2.400 ;
      LAYER via2 ;
        RECT 541.280 499.490 541.560 499.770 ;
        RECT 541.510 497.960 541.790 498.240 ;
      LAYER met3 ;
        RECT 541.255 499.620 541.585 499.795 ;
        RECT 541.230 499.610 541.610 499.620 ;
        RECT 541.230 499.310 541.870 499.610 ;
        RECT 541.230 499.300 541.610 499.310 ;
        RECT 541.485 498.260 541.815 498.265 ;
        RECT 541.230 498.250 541.815 498.260 ;
        RECT 541.030 497.950 541.815 498.250 ;
        RECT 541.230 497.940 541.815 497.950 ;
        RECT 541.485 497.935 541.815 497.940 ;
      LAYER via3 ;
        RECT 541.260 499.300 541.580 499.620 ;
        RECT 541.260 497.940 541.580 498.260 ;
      LAYER met4 ;
        RECT 541.255 499.295 541.585 499.625 ;
        RECT 541.270 498.265 541.570 499.295 ;
        RECT 541.255 497.935 541.585 498.265 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 542.640 499.700 542.960 499.760 ;
        RECT 542.500 499.500 542.960 499.700 ;
        RECT 542.500 497.380 542.640 499.500 ;
        RECT 542.410 497.120 542.730 497.380 ;
        RECT 540.110 451.080 540.430 451.140 ;
        RECT 542.870 451.080 543.190 451.140 ;
        RECT 540.110 450.940 543.190 451.080 ;
        RECT 540.110 450.880 540.430 450.940 ;
        RECT 542.870 450.880 543.190 450.940 ;
        RECT 540.110 66.880 540.430 66.940 ;
        RECT 1677.690 66.880 1678.010 66.940 ;
        RECT 540.110 66.740 1678.010 66.880 ;
        RECT 540.110 66.680 540.430 66.740 ;
        RECT 1677.690 66.680 1678.010 66.740 ;
      LAYER via ;
        RECT 542.670 499.500 542.930 499.760 ;
        RECT 542.440 497.120 542.700 497.380 ;
        RECT 540.140 450.880 540.400 451.140 ;
        RECT 542.900 450.880 543.160 451.140 ;
        RECT 540.140 66.680 540.400 66.940 ;
        RECT 1677.720 66.680 1677.980 66.940 ;
      LAYER met2 ;
        RECT 542.690 500.000 542.970 504.000 ;
        RECT 542.730 499.790 542.870 500.000 ;
        RECT 542.670 499.470 542.930 499.790 ;
        RECT 542.440 497.090 542.700 497.410 ;
        RECT 542.500 496.870 542.640 497.090 ;
        RECT 542.500 496.730 543.100 496.870 ;
        RECT 542.960 451.170 543.100 496.730 ;
        RECT 540.140 450.850 540.400 451.170 ;
        RECT 542.900 450.850 543.160 451.170 ;
        RECT 540.200 66.970 540.340 450.850 ;
        RECT 540.140 66.650 540.400 66.970 ;
        RECT 1677.720 66.650 1677.980 66.970 ;
        RECT 1677.780 2.400 1677.920 66.650 ;
        RECT 1677.570 -4.800 1678.130 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.170 500.000 468.450 504.000 ;
        RECT 468.210 499.815 468.350 500.000 ;
        RECT 468.140 499.445 468.420 499.815 ;
        RECT 783.470 58.635 783.750 59.005 ;
        RECT 783.540 2.400 783.680 58.635 ;
        RECT 783.330 -4.800 783.890 2.400 ;
      LAYER via2 ;
        RECT 468.140 499.490 468.420 499.770 ;
        RECT 783.470 58.680 783.750 58.960 ;
      LAYER met3 ;
        RECT 466.710 499.610 467.090 499.620 ;
        RECT 468.115 499.610 468.445 499.795 ;
        RECT 466.710 499.465 468.445 499.610 ;
        RECT 466.710 499.310 468.430 499.465 ;
        RECT 466.710 499.300 467.090 499.310 ;
        RECT 465.790 58.970 466.170 58.980 ;
        RECT 783.445 58.970 783.775 58.985 ;
        RECT 465.790 58.670 783.775 58.970 ;
        RECT 465.790 58.660 466.170 58.670 ;
        RECT 783.445 58.655 783.775 58.670 ;
      LAYER via3 ;
        RECT 466.740 499.300 467.060 499.620 ;
        RECT 465.820 58.660 466.140 58.980 ;
      LAYER met4 ;
        RECT 466.735 499.610 467.065 499.625 ;
        RECT 465.830 499.310 467.065 499.610 ;
        RECT 465.830 58.985 466.130 499.310 ;
        RECT 466.735 499.295 467.065 499.310 ;
        RECT 465.815 58.655 466.145 58.985 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.070 500.000 544.350 504.000 ;
        RECT 544.110 499.475 544.250 500.000 ;
        RECT 544.040 499.105 544.320 499.475 ;
        RECT 543.810 497.235 544.090 497.605 ;
        RECT 543.880 483.325 544.020 497.235 ;
        RECT 543.810 482.955 544.090 483.325 ;
        RECT 1694.270 65.435 1694.550 65.805 ;
        RECT 1694.340 2.400 1694.480 65.435 ;
        RECT 1694.130 -4.800 1694.690 2.400 ;
      LAYER via2 ;
        RECT 544.040 499.150 544.320 499.430 ;
        RECT 543.810 497.280 544.090 497.560 ;
        RECT 543.810 483.000 544.090 483.280 ;
        RECT 1694.270 65.480 1694.550 65.760 ;
      LAYER met3 ;
        RECT 544.015 499.125 544.345 499.455 ;
        RECT 544.030 497.585 544.330 499.125 ;
        RECT 543.785 497.270 544.330 497.585 ;
        RECT 543.785 497.255 544.115 497.270 ;
        RECT 543.785 483.300 544.115 483.305 ;
        RECT 543.785 483.290 544.370 483.300 ;
        RECT 543.785 482.990 544.570 483.290 ;
        RECT 543.785 482.980 544.370 482.990 ;
        RECT 543.785 482.975 544.115 482.980 ;
        RECT 543.990 65.770 544.370 65.780 ;
        RECT 1694.245 65.770 1694.575 65.785 ;
        RECT 543.990 65.470 1694.575 65.770 ;
        RECT 543.990 65.460 544.370 65.470 ;
        RECT 1694.245 65.455 1694.575 65.470 ;
      LAYER via3 ;
        RECT 544.020 482.980 544.340 483.300 ;
        RECT 544.020 65.460 544.340 65.780 ;
      LAYER met4 ;
        RECT 544.015 482.975 544.345 483.305 ;
        RECT 544.030 65.785 544.330 482.975 ;
        RECT 544.015 65.455 544.345 65.785 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.400 499.500 545.720 499.760 ;
        RECT 545.490 498.400 545.630 499.500 ;
        RECT 545.170 498.200 545.630 498.400 ;
        RECT 545.170 498.140 545.490 498.200 ;
        RECT 545.170 480.660 545.490 480.720 ;
        RECT 547.470 480.660 547.790 480.720 ;
        RECT 545.170 480.520 547.790 480.660 ;
        RECT 545.170 480.460 545.490 480.520 ;
        RECT 547.470 480.460 547.790 480.520 ;
        RECT 547.470 156.300 547.790 156.360 ;
        RECT 1704.830 156.300 1705.150 156.360 ;
        RECT 547.470 156.160 1705.150 156.300 ;
        RECT 547.470 156.100 547.790 156.160 ;
        RECT 1704.830 156.100 1705.150 156.160 ;
        RECT 1704.830 20.300 1705.150 20.360 ;
        RECT 1710.810 20.300 1711.130 20.360 ;
        RECT 1704.830 20.160 1711.130 20.300 ;
        RECT 1704.830 20.100 1705.150 20.160 ;
        RECT 1710.810 20.100 1711.130 20.160 ;
      LAYER via ;
        RECT 545.430 499.500 545.690 499.760 ;
        RECT 545.200 498.140 545.460 498.400 ;
        RECT 545.200 480.460 545.460 480.720 ;
        RECT 547.500 480.460 547.760 480.720 ;
        RECT 547.500 156.100 547.760 156.360 ;
        RECT 1704.860 156.100 1705.120 156.360 ;
        RECT 1704.860 20.100 1705.120 20.360 ;
        RECT 1710.840 20.100 1711.100 20.360 ;
      LAYER met2 ;
        RECT 545.450 500.000 545.730 504.000 ;
        RECT 545.490 499.790 545.630 500.000 ;
        RECT 545.430 499.470 545.690 499.790 ;
        RECT 545.200 498.110 545.460 498.430 ;
        RECT 545.260 480.750 545.400 498.110 ;
        RECT 545.200 480.430 545.460 480.750 ;
        RECT 547.500 480.430 547.760 480.750 ;
        RECT 547.560 156.390 547.700 480.430 ;
        RECT 547.500 156.070 547.760 156.390 ;
        RECT 1704.860 156.070 1705.120 156.390 ;
        RECT 1704.920 20.390 1705.060 156.070 ;
        RECT 1704.860 20.070 1705.120 20.390 ;
        RECT 1710.840 20.070 1711.100 20.390 ;
        RECT 1710.900 2.400 1711.040 20.070 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.780 499.160 547.100 499.420 ;
        RECT 546.870 497.320 547.010 499.160 ;
        RECT 548.390 497.320 548.710 497.380 ;
        RECT 546.870 497.180 548.710 497.320 ;
        RECT 548.390 497.120 548.710 497.180 ;
        RECT 548.390 417.420 548.710 417.480 ;
        RECT 1725.070 417.420 1725.390 417.480 ;
        RECT 548.390 417.280 1725.390 417.420 ;
        RECT 548.390 417.220 548.710 417.280 ;
        RECT 1725.070 417.220 1725.390 417.280 ;
      LAYER via ;
        RECT 546.810 499.160 547.070 499.420 ;
        RECT 548.420 497.120 548.680 497.380 ;
        RECT 548.420 417.220 548.680 417.480 ;
        RECT 1725.100 417.220 1725.360 417.480 ;
      LAYER met2 ;
        RECT 546.830 500.000 547.110 504.000 ;
        RECT 546.870 499.450 547.010 500.000 ;
        RECT 546.810 499.130 547.070 499.450 ;
        RECT 548.420 497.090 548.680 497.410 ;
        RECT 548.480 417.510 548.620 497.090 ;
        RECT 548.420 417.190 548.680 417.510 ;
        RECT 1725.100 417.190 1725.360 417.510 ;
        RECT 1725.160 82.870 1725.300 417.190 ;
        RECT 1725.160 82.730 1727.600 82.870 ;
        RECT 1727.460 2.400 1727.600 82.730 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 547.930 472.840 548.250 472.900 ;
        RECT 544.800 472.700 548.250 472.840 ;
        RECT 544.800 472.560 544.940 472.700 ;
        RECT 547.930 472.640 548.250 472.700 ;
        RECT 544.710 472.300 545.030 472.560 ;
        RECT 545.170 59.060 545.490 59.120 ;
        RECT 1743.930 59.060 1744.250 59.120 ;
        RECT 545.170 58.920 1744.250 59.060 ;
        RECT 545.170 58.860 545.490 58.920 ;
        RECT 1743.930 58.860 1744.250 58.920 ;
      LAYER via ;
        RECT 547.960 472.640 548.220 472.900 ;
        RECT 544.740 472.300 545.000 472.560 ;
        RECT 545.200 58.860 545.460 59.120 ;
        RECT 1743.960 58.860 1744.220 59.120 ;
      LAYER met2 ;
        RECT 548.210 500.000 548.490 504.000 ;
        RECT 548.250 498.680 548.390 500.000 ;
        RECT 548.020 498.540 548.390 498.680 ;
        RECT 548.020 472.930 548.160 498.540 ;
        RECT 547.960 472.610 548.220 472.930 ;
        RECT 544.740 472.270 545.000 472.590 ;
        RECT 544.800 462.370 544.940 472.270 ;
        RECT 544.800 462.230 545.400 462.370 ;
        RECT 545.260 59.150 545.400 462.230 ;
        RECT 545.200 58.830 545.460 59.150 ;
        RECT 1743.960 58.830 1744.220 59.150 ;
        RECT 1744.020 2.400 1744.160 58.830 ;
        RECT 1743.810 -4.800 1744.370 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.540 500.040 549.860 500.100 ;
        RECT 548.710 499.900 549.860 500.040 ;
        RECT 548.710 497.660 548.850 499.900 ;
        RECT 549.540 499.840 549.860 499.900 ;
        RECT 549.770 497.660 550.090 497.720 ;
        RECT 548.710 497.520 550.090 497.660 ;
        RECT 549.770 497.460 550.090 497.520 ;
        RECT 547.010 478.280 547.330 478.340 ;
        RECT 549.770 478.280 550.090 478.340 ;
        RECT 547.010 478.140 550.090 478.280 ;
        RECT 547.010 478.080 547.330 478.140 ;
        RECT 549.770 478.080 550.090 478.140 ;
        RECT 547.010 74.020 547.330 74.080 ;
        RECT 1760.490 74.020 1760.810 74.080 ;
        RECT 547.010 73.880 1760.810 74.020 ;
        RECT 547.010 73.820 547.330 73.880 ;
        RECT 1760.490 73.820 1760.810 73.880 ;
      LAYER via ;
        RECT 549.570 499.840 549.830 500.100 ;
        RECT 549.800 497.460 550.060 497.720 ;
        RECT 547.040 478.080 547.300 478.340 ;
        RECT 549.800 478.080 550.060 478.340 ;
        RECT 547.040 73.820 547.300 74.080 ;
        RECT 1760.520 73.820 1760.780 74.080 ;
      LAYER met2 ;
        RECT 549.590 500.130 549.870 504.000 ;
        RECT 549.570 500.000 549.870 500.130 ;
        RECT 549.570 499.810 549.830 500.000 ;
        RECT 549.800 497.430 550.060 497.750 ;
        RECT 549.860 478.370 550.000 497.430 ;
        RECT 547.040 478.050 547.300 478.370 ;
        RECT 549.800 478.050 550.060 478.370 ;
        RECT 547.100 74.110 547.240 478.050 ;
        RECT 547.040 73.790 547.300 74.110 ;
        RECT 1760.520 73.790 1760.780 74.110 ;
        RECT 1760.580 2.400 1760.720 73.790 ;
        RECT 1760.370 -4.800 1760.930 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 551.610 468.760 551.930 468.820 ;
        RECT 557.590 468.760 557.910 468.820 ;
        RECT 551.610 468.620 557.910 468.760 ;
        RECT 551.610 468.560 551.930 468.620 ;
        RECT 557.590 468.560 557.910 468.620 ;
        RECT 557.130 155.960 557.450 156.020 ;
        RECT 1773.370 155.960 1773.690 156.020 ;
        RECT 557.130 155.820 1773.690 155.960 ;
        RECT 557.130 155.760 557.450 155.820 ;
        RECT 1773.370 155.760 1773.690 155.820 ;
      LAYER via ;
        RECT 551.640 468.560 551.900 468.820 ;
        RECT 557.620 468.560 557.880 468.820 ;
        RECT 557.160 155.760 557.420 156.020 ;
        RECT 1773.400 155.760 1773.660 156.020 ;
      LAYER met2 ;
        RECT 550.970 500.000 551.250 504.000 ;
        RECT 551.010 499.645 551.150 500.000 ;
        RECT 550.940 499.275 551.220 499.645 ;
        RECT 551.630 490.435 551.910 490.805 ;
        RECT 551.700 468.850 551.840 490.435 ;
        RECT 551.640 468.530 551.900 468.850 ;
        RECT 557.620 468.530 557.880 468.850 ;
        RECT 557.680 420.970 557.820 468.530 ;
        RECT 557.220 420.830 557.820 420.970 ;
        RECT 557.220 156.050 557.360 420.830 ;
        RECT 557.160 155.730 557.420 156.050 ;
        RECT 1773.400 155.730 1773.660 156.050 ;
        RECT 1773.460 82.870 1773.600 155.730 ;
        RECT 1773.460 82.730 1777.280 82.870 ;
        RECT 1777.140 2.400 1777.280 82.730 ;
        RECT 1776.930 -4.800 1777.490 2.400 ;
      LAYER via2 ;
        RECT 550.940 499.320 551.220 499.600 ;
        RECT 551.630 490.480 551.910 490.760 ;
      LAYER met3 ;
        RECT 549.510 499.610 549.890 499.620 ;
        RECT 550.915 499.610 551.245 499.625 ;
        RECT 549.510 499.310 551.245 499.610 ;
        RECT 549.510 499.300 549.890 499.310 ;
        RECT 550.915 499.295 551.245 499.310 ;
        RECT 550.430 490.770 550.810 490.780 ;
        RECT 551.605 490.770 551.935 490.785 ;
        RECT 550.430 490.470 551.935 490.770 ;
        RECT 550.430 490.460 550.810 490.470 ;
        RECT 551.605 490.455 551.935 490.470 ;
      LAYER via3 ;
        RECT 549.540 499.300 549.860 499.620 ;
        RECT 550.460 490.460 550.780 490.780 ;
      LAYER met4 ;
        RECT 549.535 499.610 549.865 499.625 ;
        RECT 549.535 499.310 550.770 499.610 ;
        RECT 549.535 499.295 549.865 499.310 ;
        RECT 550.470 490.785 550.770 499.310 ;
        RECT 550.455 490.455 550.785 490.785 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.300 499.700 552.620 499.760 ;
        RECT 552.300 499.560 553.680 499.700 ;
        RECT 552.300 499.500 552.620 499.560 ;
        RECT 553.540 497.720 553.680 499.560 ;
        RECT 553.450 497.460 553.770 497.720 ;
        RECT 553.450 141.340 553.770 141.400 ;
        RECT 1787.630 141.340 1787.950 141.400 ;
        RECT 553.450 141.200 1787.950 141.340 ;
        RECT 553.450 141.140 553.770 141.200 ;
        RECT 1787.630 141.140 1787.950 141.200 ;
        RECT 1787.630 20.300 1787.950 20.360 ;
        RECT 1793.610 20.300 1793.930 20.360 ;
        RECT 1787.630 20.160 1793.930 20.300 ;
        RECT 1787.630 20.100 1787.950 20.160 ;
        RECT 1793.610 20.100 1793.930 20.160 ;
      LAYER via ;
        RECT 552.330 499.500 552.590 499.760 ;
        RECT 553.480 497.460 553.740 497.720 ;
        RECT 553.480 141.140 553.740 141.400 ;
        RECT 1787.660 141.140 1787.920 141.400 ;
        RECT 1787.660 20.100 1787.920 20.360 ;
        RECT 1793.640 20.100 1793.900 20.360 ;
      LAYER met2 ;
        RECT 552.350 500.000 552.630 504.000 ;
        RECT 552.390 499.790 552.530 500.000 ;
        RECT 552.330 499.470 552.590 499.790 ;
        RECT 553.480 497.430 553.740 497.750 ;
        RECT 553.540 141.430 553.680 497.430 ;
        RECT 553.480 141.110 553.740 141.430 ;
        RECT 1787.660 141.110 1787.920 141.430 ;
        RECT 1787.720 20.390 1787.860 141.110 ;
        RECT 1787.660 20.070 1787.920 20.390 ;
        RECT 1793.640 20.070 1793.900 20.390 ;
        RECT 1793.700 2.400 1793.840 20.070 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.910 155.620 554.230 155.680 ;
        RECT 1807.870 155.620 1808.190 155.680 ;
        RECT 553.910 155.480 1808.190 155.620 ;
        RECT 553.910 155.420 554.230 155.480 ;
        RECT 1807.870 155.420 1808.190 155.480 ;
      LAYER via ;
        RECT 553.940 155.420 554.200 155.680 ;
        RECT 1807.900 155.420 1808.160 155.680 ;
      LAYER met2 ;
        RECT 553.730 500.000 554.010 504.000 ;
        RECT 553.770 499.020 553.910 500.000 ;
        RECT 553.770 498.880 554.140 499.020 ;
        RECT 554.000 155.710 554.140 498.880 ;
        RECT 553.940 155.390 554.200 155.710 ;
        RECT 1807.900 155.390 1808.160 155.710 ;
        RECT 1807.960 82.870 1808.100 155.390 ;
        RECT 1807.960 82.730 1810.400 82.870 ;
        RECT 1810.260 2.400 1810.400 82.730 ;
        RECT 1810.050 -4.800 1810.610 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.060 499.500 555.380 499.760 ;
        RECT 555.150 498.340 555.290 499.500 ;
        RECT 555.150 498.200 555.980 498.340 ;
        RECT 554.370 497.660 554.690 497.720 ;
        RECT 555.840 497.660 555.980 498.200 ;
        RECT 554.370 497.520 555.980 497.660 ;
        RECT 554.370 497.460 554.690 497.520 ;
        RECT 554.370 155.280 554.690 155.340 ;
        RECT 1821.670 155.280 1821.990 155.340 ;
        RECT 554.370 155.140 1821.990 155.280 ;
        RECT 554.370 155.080 554.690 155.140 ;
        RECT 1821.670 155.080 1821.990 155.140 ;
      LAYER via ;
        RECT 555.090 499.500 555.350 499.760 ;
        RECT 554.400 497.460 554.660 497.720 ;
        RECT 554.400 155.080 554.660 155.340 ;
        RECT 1821.700 155.080 1821.960 155.340 ;
      LAYER met2 ;
        RECT 555.110 500.000 555.390 504.000 ;
        RECT 555.150 499.790 555.290 500.000 ;
        RECT 555.090 499.470 555.350 499.790 ;
        RECT 554.400 497.430 554.660 497.750 ;
        RECT 554.460 155.370 554.600 497.430 ;
        RECT 554.400 155.050 554.660 155.370 ;
        RECT 1821.700 155.050 1821.960 155.370 ;
        RECT 1821.760 82.870 1821.900 155.050 ;
        RECT 1821.760 82.730 1826.960 82.870 ;
        RECT 1826.820 2.400 1826.960 82.730 ;
        RECT 1826.610 -4.800 1827.170 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 556.670 498.000 556.990 498.060 ;
        RECT 557.590 498.000 557.910 498.060 ;
        RECT 556.670 497.860 557.910 498.000 ;
        RECT 556.670 497.800 556.990 497.860 ;
        RECT 557.590 497.800 557.910 497.860 ;
        RECT 552.530 477.940 552.850 478.000 ;
        RECT 557.590 477.940 557.910 478.000 ;
        RECT 552.530 477.800 557.910 477.940 ;
        RECT 552.530 477.740 552.850 477.800 ;
        RECT 557.590 477.740 557.910 477.800 ;
        RECT 552.530 73.680 552.850 73.740 ;
        RECT 1843.290 73.680 1843.610 73.740 ;
        RECT 552.530 73.540 1843.610 73.680 ;
        RECT 552.530 73.480 552.850 73.540 ;
        RECT 1843.290 73.480 1843.610 73.540 ;
      LAYER via ;
        RECT 556.700 497.800 556.960 498.060 ;
        RECT 557.620 497.800 557.880 498.060 ;
        RECT 552.560 477.740 552.820 478.000 ;
        RECT 557.620 477.740 557.880 478.000 ;
        RECT 552.560 73.480 552.820 73.740 ;
        RECT 1843.320 73.480 1843.580 73.740 ;
      LAYER met2 ;
        RECT 556.490 500.000 556.770 504.000 ;
        RECT 556.530 498.850 556.670 500.000 ;
        RECT 556.530 498.710 556.900 498.850 ;
        RECT 556.760 498.090 556.900 498.710 ;
        RECT 556.700 497.770 556.960 498.090 ;
        RECT 557.620 497.770 557.880 498.090 ;
        RECT 557.680 478.030 557.820 497.770 ;
        RECT 552.560 477.710 552.820 478.030 ;
        RECT 557.620 477.710 557.880 478.030 ;
        RECT 552.620 73.770 552.760 477.710 ;
        RECT 552.560 73.450 552.820 73.770 ;
        RECT 1843.320 73.450 1843.580 73.770 ;
        RECT 1843.380 2.400 1843.520 73.450 ;
        RECT 1843.170 -4.800 1843.730 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.500 499.500 469.820 499.760 ;
        RECT 469.590 498.400 469.730 499.500 ;
        RECT 469.270 498.200 469.730 498.400 ;
        RECT 469.270 498.140 469.590 498.200 ;
        RECT 468.810 472.160 469.130 472.220 ;
        RECT 470.190 472.160 470.510 472.220 ;
        RECT 468.810 472.020 470.510 472.160 ;
        RECT 468.810 471.960 469.130 472.020 ;
        RECT 470.190 471.960 470.510 472.020 ;
        RECT 470.190 157.660 470.510 157.720 ;
        RECT 794.030 157.660 794.350 157.720 ;
        RECT 470.190 157.520 794.350 157.660 ;
        RECT 470.190 157.460 470.510 157.520 ;
        RECT 794.030 157.460 794.350 157.520 ;
        RECT 794.030 19.960 794.350 20.020 ;
        RECT 800.010 19.960 800.330 20.020 ;
        RECT 794.030 19.820 800.330 19.960 ;
        RECT 794.030 19.760 794.350 19.820 ;
        RECT 800.010 19.760 800.330 19.820 ;
      LAYER via ;
        RECT 469.530 499.500 469.790 499.760 ;
        RECT 469.300 498.140 469.560 498.400 ;
        RECT 468.840 471.960 469.100 472.220 ;
        RECT 470.220 471.960 470.480 472.220 ;
        RECT 470.220 157.460 470.480 157.720 ;
        RECT 794.060 157.460 794.320 157.720 ;
        RECT 794.060 19.760 794.320 20.020 ;
        RECT 800.040 19.760 800.300 20.020 ;
      LAYER met2 ;
        RECT 469.550 500.000 469.830 504.000 ;
        RECT 469.590 499.790 469.730 500.000 ;
        RECT 469.530 499.470 469.790 499.790 ;
        RECT 469.300 498.110 469.560 498.430 ;
        RECT 469.360 473.690 469.500 498.110 ;
        RECT 468.900 473.550 469.500 473.690 ;
        RECT 468.900 472.250 469.040 473.550 ;
        RECT 468.840 471.930 469.100 472.250 ;
        RECT 470.220 471.930 470.480 472.250 ;
        RECT 470.280 157.750 470.420 471.930 ;
        RECT 470.220 157.430 470.480 157.750 ;
        RECT 794.060 157.430 794.320 157.750 ;
        RECT 794.120 20.050 794.260 157.430 ;
        RECT 794.060 19.730 794.320 20.050 ;
        RECT 800.040 19.730 800.300 20.050 ;
        RECT 800.100 2.400 800.240 19.730 ;
        RECT 799.890 -4.800 800.450 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 557.820 499.700 558.140 499.760 ;
        RECT 557.820 499.560 558.970 499.700 ;
        RECT 557.820 499.500 558.140 499.560 ;
        RECT 558.830 498.060 558.970 499.560 ;
        RECT 558.510 497.860 558.970 498.060 ;
        RECT 558.510 497.800 558.830 497.860 ;
      LAYER via ;
        RECT 557.850 499.500 558.110 499.760 ;
        RECT 558.540 497.800 558.800 498.060 ;
      LAYER met2 ;
        RECT 557.870 500.000 558.150 504.000 ;
        RECT 557.910 499.790 558.050 500.000 ;
        RECT 557.850 499.470 558.110 499.790 ;
        RECT 558.540 497.770 558.800 498.090 ;
        RECT 558.600 481.965 558.740 497.770 ;
        RECT 558.530 481.595 558.810 481.965 ;
        RECT 1859.870 73.595 1860.150 73.965 ;
        RECT 1859.940 2.400 1860.080 73.595 ;
        RECT 1859.730 -4.800 1860.290 2.400 ;
      LAYER via2 ;
        RECT 558.530 481.640 558.810 481.920 ;
        RECT 1859.870 73.640 1860.150 73.920 ;
      LAYER met3 ;
        RECT 555.030 481.930 555.410 481.940 ;
        RECT 558.505 481.930 558.835 481.945 ;
        RECT 555.030 481.630 558.835 481.930 ;
        RECT 555.030 481.620 555.410 481.630 ;
        RECT 558.505 481.615 558.835 481.630 ;
        RECT 555.030 73.930 555.410 73.940 ;
        RECT 1859.845 73.930 1860.175 73.945 ;
        RECT 555.030 73.630 1860.175 73.930 ;
        RECT 555.030 73.620 555.410 73.630 ;
        RECT 1859.845 73.615 1860.175 73.630 ;
      LAYER via3 ;
        RECT 555.060 481.620 555.380 481.940 ;
        RECT 555.060 73.620 555.380 73.940 ;
      LAYER met4 ;
        RECT 555.055 481.615 555.385 481.945 ;
        RECT 555.070 73.945 555.370 481.615 ;
        RECT 555.055 73.615 555.385 73.945 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.200 499.160 559.520 499.420 ;
        RECT 558.050 496.300 558.370 496.360 ;
        RECT 559.290 496.300 559.430 499.160 ;
        RECT 558.050 496.160 559.430 496.300 ;
        RECT 558.050 496.100 558.370 496.160 ;
        RECT 558.050 484.060 558.370 484.120 ;
        RECT 564.030 484.060 564.350 484.120 ;
        RECT 558.050 483.920 564.350 484.060 ;
        RECT 558.050 483.860 558.370 483.920 ;
        RECT 564.030 483.860 564.350 483.920 ;
        RECT 564.030 466.380 564.350 466.440 ;
        RECT 1869.970 466.380 1870.290 466.440 ;
        RECT 564.030 466.240 1870.290 466.380 ;
        RECT 564.030 466.180 564.350 466.240 ;
        RECT 1869.970 466.180 1870.290 466.240 ;
        RECT 1869.970 16.900 1870.290 16.960 ;
        RECT 1876.410 16.900 1876.730 16.960 ;
        RECT 1869.970 16.760 1876.730 16.900 ;
        RECT 1869.970 16.700 1870.290 16.760 ;
        RECT 1876.410 16.700 1876.730 16.760 ;
      LAYER via ;
        RECT 559.230 499.160 559.490 499.420 ;
        RECT 558.080 496.100 558.340 496.360 ;
        RECT 558.080 483.860 558.340 484.120 ;
        RECT 564.060 483.860 564.320 484.120 ;
        RECT 564.060 466.180 564.320 466.440 ;
        RECT 1870.000 466.180 1870.260 466.440 ;
        RECT 1870.000 16.700 1870.260 16.960 ;
        RECT 1876.440 16.700 1876.700 16.960 ;
      LAYER met2 ;
        RECT 559.250 500.000 559.530 504.000 ;
        RECT 559.290 499.450 559.430 500.000 ;
        RECT 559.230 499.130 559.490 499.450 ;
        RECT 558.080 496.070 558.340 496.390 ;
        RECT 558.140 484.150 558.280 496.070 ;
        RECT 558.080 483.830 558.340 484.150 ;
        RECT 564.060 483.830 564.320 484.150 ;
        RECT 564.120 466.470 564.260 483.830 ;
        RECT 564.060 466.150 564.320 466.470 ;
        RECT 1870.000 466.150 1870.260 466.470 ;
        RECT 1870.060 16.990 1870.200 466.150 ;
        RECT 1870.000 16.670 1870.260 16.990 ;
        RECT 1876.440 16.670 1876.700 16.990 ;
        RECT 1876.500 2.400 1876.640 16.670 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.270 163.780 561.590 163.840 ;
        RECT 1890.670 163.780 1890.990 163.840 ;
        RECT 561.270 163.640 1890.990 163.780 ;
        RECT 561.270 163.580 561.590 163.640 ;
        RECT 1890.670 163.580 1890.990 163.640 ;
      LAYER via ;
        RECT 561.300 163.580 561.560 163.840 ;
        RECT 1890.700 163.580 1890.960 163.840 ;
      LAYER met2 ;
        RECT 560.630 500.000 560.910 504.000 ;
        RECT 560.670 498.850 560.810 500.000 ;
        RECT 560.440 498.710 560.810 498.850 ;
        RECT 560.440 498.285 560.580 498.710 ;
        RECT 560.370 497.915 560.650 498.285 ;
        RECT 561.290 496.555 561.570 496.925 ;
        RECT 561.360 163.870 561.500 496.555 ;
        RECT 561.300 163.550 561.560 163.870 ;
        RECT 1890.700 163.550 1890.960 163.870 ;
        RECT 1890.760 82.870 1890.900 163.550 ;
        RECT 1890.760 82.730 1893.200 82.870 ;
        RECT 1893.060 2.400 1893.200 82.730 ;
        RECT 1892.850 -4.800 1893.410 2.400 ;
      LAYER via2 ;
        RECT 560.370 497.960 560.650 498.240 ;
        RECT 561.290 496.600 561.570 496.880 ;
      LAYER met3 ;
        RECT 560.345 498.250 560.675 498.265 ;
        RECT 560.345 497.935 560.890 498.250 ;
        RECT 560.590 496.890 560.890 497.935 ;
        RECT 561.265 496.890 561.595 496.905 ;
        RECT 560.590 496.590 561.595 496.890 ;
        RECT 561.265 496.575 561.595 496.590 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 561.730 163.440 562.050 163.500 ;
        RECT 1904.470 163.440 1904.790 163.500 ;
        RECT 561.730 163.300 1904.790 163.440 ;
        RECT 561.730 163.240 562.050 163.300 ;
        RECT 1904.470 163.240 1904.790 163.300 ;
      LAYER via ;
        RECT 561.760 163.240 562.020 163.500 ;
        RECT 1904.500 163.240 1904.760 163.500 ;
      LAYER met2 ;
        RECT 562.010 500.000 562.290 504.000 ;
        RECT 562.050 498.850 562.190 500.000 ;
        RECT 561.820 498.710 562.190 498.850 ;
        RECT 561.820 163.530 561.960 498.710 ;
        RECT 561.760 163.210 562.020 163.530 ;
        RECT 1904.500 163.210 1904.760 163.530 ;
        RECT 1904.560 82.870 1904.700 163.210 ;
        RECT 1904.560 82.730 1909.760 82.870 ;
        RECT 1909.620 2.400 1909.760 82.730 ;
        RECT 1909.410 -4.800 1909.970 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.810 471.820 561.130 471.880 ;
        RECT 562.650 471.820 562.970 471.880 ;
        RECT 560.810 471.680 562.970 471.820 ;
        RECT 560.810 471.620 561.130 471.680 ;
        RECT 562.650 471.620 562.970 471.680 ;
        RECT 560.810 163.100 561.130 163.160 ;
        RECT 1925.630 163.100 1925.950 163.160 ;
        RECT 560.810 162.960 1925.950 163.100 ;
        RECT 560.810 162.900 561.130 162.960 ;
        RECT 1925.630 162.900 1925.950 162.960 ;
      LAYER via ;
        RECT 560.840 471.620 561.100 471.880 ;
        RECT 562.680 471.620 562.940 471.880 ;
        RECT 560.840 162.900 561.100 163.160 ;
        RECT 1925.660 162.900 1925.920 163.160 ;
      LAYER met2 ;
        RECT 563.390 500.000 563.670 504.000 ;
        RECT 563.430 499.530 563.570 500.000 ;
        RECT 563.200 499.390 563.570 499.530 ;
        RECT 563.200 497.490 563.340 499.390 ;
        RECT 562.740 497.350 563.340 497.490 ;
        RECT 562.740 471.910 562.880 497.350 ;
        RECT 560.840 471.590 561.100 471.910 ;
        RECT 562.680 471.590 562.940 471.910 ;
        RECT 560.900 163.190 561.040 471.590 ;
        RECT 560.840 162.870 561.100 163.190 ;
        RECT 1925.660 162.870 1925.920 163.190 ;
        RECT 1925.720 82.870 1925.860 162.870 ;
        RECT 1925.720 82.730 1926.320 82.870 ;
        RECT 1926.180 2.400 1926.320 82.730 ;
        RECT 1925.970 -4.800 1926.530 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.770 500.000 565.050 504.000 ;
        RECT 564.810 498.340 564.950 500.000 ;
        RECT 564.810 498.200 565.180 498.340 ;
        RECT 565.040 497.490 565.180 498.200 ;
        RECT 564.580 497.350 565.180 497.490 ;
        RECT 564.580 483.325 564.720 497.350 ;
        RECT 564.510 482.955 564.790 483.325 ;
        RECT 1942.670 72.235 1942.950 72.605 ;
        RECT 1942.740 2.400 1942.880 72.235 ;
        RECT 1942.530 -4.800 1943.090 2.400 ;
      LAYER via2 ;
        RECT 564.510 483.000 564.790 483.280 ;
        RECT 1942.670 72.280 1942.950 72.560 ;
      LAYER met3 ;
        RECT 564.485 483.300 564.815 483.305 ;
        RECT 564.230 483.290 564.815 483.300 ;
        RECT 564.030 482.990 564.815 483.290 ;
        RECT 564.230 482.980 564.815 482.990 ;
        RECT 564.485 482.975 564.815 482.980 ;
        RECT 564.230 72.570 564.610 72.580 ;
        RECT 1942.645 72.570 1942.975 72.585 ;
        RECT 564.230 72.270 1942.975 72.570 ;
        RECT 564.230 72.260 564.610 72.270 ;
        RECT 1942.645 72.255 1942.975 72.270 ;
      LAYER via3 ;
        RECT 564.260 482.980 564.580 483.300 ;
        RECT 564.260 72.260 564.580 72.580 ;
      LAYER met4 ;
        RECT 564.255 482.975 564.585 483.305 ;
        RECT 564.270 72.585 564.570 482.975 ;
        RECT 564.255 72.255 564.585 72.585 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.410 471.820 565.730 471.880 ;
        RECT 568.630 471.820 568.950 471.880 ;
        RECT 565.410 471.680 568.950 471.820 ;
        RECT 565.410 471.620 565.730 471.680 ;
        RECT 568.630 471.620 568.950 471.680 ;
        RECT 568.630 162.760 568.950 162.820 ;
        RECT 1953.230 162.760 1953.550 162.820 ;
        RECT 568.630 162.620 1953.550 162.760 ;
        RECT 568.630 162.560 568.950 162.620 ;
        RECT 1953.230 162.560 1953.550 162.620 ;
        RECT 1953.230 20.300 1953.550 20.360 ;
        RECT 1959.210 20.300 1959.530 20.360 ;
        RECT 1953.230 20.160 1959.530 20.300 ;
        RECT 1953.230 20.100 1953.550 20.160 ;
        RECT 1959.210 20.100 1959.530 20.160 ;
      LAYER via ;
        RECT 565.440 471.620 565.700 471.880 ;
        RECT 568.660 471.620 568.920 471.880 ;
        RECT 568.660 162.560 568.920 162.820 ;
        RECT 1953.260 162.560 1953.520 162.820 ;
        RECT 1953.260 20.100 1953.520 20.360 ;
        RECT 1959.240 20.100 1959.500 20.360 ;
      LAYER met2 ;
        RECT 566.150 500.000 566.430 504.000 ;
        RECT 566.190 498.850 566.330 500.000 ;
        RECT 565.960 498.710 566.330 498.850 ;
        RECT 565.960 473.690 566.100 498.710 ;
        RECT 565.500 473.550 566.100 473.690 ;
        RECT 565.500 471.910 565.640 473.550 ;
        RECT 565.440 471.590 565.700 471.910 ;
        RECT 568.660 471.590 568.920 471.910 ;
        RECT 568.720 162.850 568.860 471.590 ;
        RECT 568.660 162.530 568.920 162.850 ;
        RECT 1953.260 162.530 1953.520 162.850 ;
        RECT 1953.320 20.390 1953.460 162.530 ;
        RECT 1953.260 20.070 1953.520 20.390 ;
        RECT 1959.240 20.070 1959.500 20.390 ;
        RECT 1959.300 2.400 1959.440 20.070 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.480 499.160 567.800 499.420 ;
        RECT 567.570 498.340 567.710 499.160 ;
        RECT 568.170 498.340 568.490 498.400 ;
        RECT 567.570 498.200 568.490 498.340 ;
        RECT 568.170 498.140 568.490 498.200 ;
        RECT 568.170 162.420 568.490 162.480 ;
        RECT 1973.470 162.420 1973.790 162.480 ;
        RECT 568.170 162.280 1973.790 162.420 ;
        RECT 568.170 162.220 568.490 162.280 ;
        RECT 1973.470 162.220 1973.790 162.280 ;
      LAYER via ;
        RECT 567.510 499.160 567.770 499.420 ;
        RECT 568.200 498.140 568.460 498.400 ;
        RECT 568.200 162.220 568.460 162.480 ;
        RECT 1973.500 162.220 1973.760 162.480 ;
      LAYER met2 ;
        RECT 567.530 500.000 567.810 504.000 ;
        RECT 567.570 499.450 567.710 500.000 ;
        RECT 567.510 499.130 567.770 499.450 ;
        RECT 568.200 498.110 568.460 498.430 ;
        RECT 568.260 162.510 568.400 498.110 ;
        RECT 568.200 162.190 568.460 162.510 ;
        RECT 1973.500 162.190 1973.760 162.510 ;
        RECT 1973.560 82.870 1973.700 162.190 ;
        RECT 1973.560 82.730 1976.000 82.870 ;
        RECT 1975.860 2.400 1976.000 82.730 ;
        RECT 1975.650 -4.800 1976.210 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.710 472.500 568.030 472.560 ;
        RECT 568.630 472.500 568.950 472.560 ;
        RECT 567.710 472.360 568.950 472.500 ;
        RECT 567.710 472.300 568.030 472.360 ;
        RECT 568.630 472.300 568.950 472.360 ;
        RECT 567.710 162.080 568.030 162.140 ;
        RECT 1987.270 162.080 1987.590 162.140 ;
        RECT 567.710 161.940 1987.590 162.080 ;
        RECT 567.710 161.880 568.030 161.940 ;
        RECT 1987.270 161.880 1987.590 161.940 ;
      LAYER via ;
        RECT 567.740 472.300 568.000 472.560 ;
        RECT 568.660 472.300 568.920 472.560 ;
        RECT 567.740 161.880 568.000 162.140 ;
        RECT 1987.300 161.880 1987.560 162.140 ;
      LAYER met2 ;
        RECT 568.910 500.000 569.190 504.000 ;
        RECT 568.950 498.850 569.090 500.000 ;
        RECT 568.720 498.710 569.090 498.850 ;
        RECT 568.720 472.590 568.860 498.710 ;
        RECT 567.740 472.270 568.000 472.590 ;
        RECT 568.660 472.270 568.920 472.590 ;
        RECT 567.800 162.170 567.940 472.270 ;
        RECT 567.740 161.850 568.000 162.170 ;
        RECT 1987.300 161.850 1987.560 162.170 ;
        RECT 1987.360 82.870 1987.500 161.850 ;
        RECT 1987.360 82.730 1992.560 82.870 ;
        RECT 1992.420 2.400 1992.560 82.730 ;
        RECT 1992.210 -4.800 1992.770 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.290 500.000 570.570 504.000 ;
        RECT 570.330 498.850 570.470 500.000 ;
        RECT 570.100 498.710 570.470 498.850 ;
        RECT 570.100 483.325 570.240 498.710 ;
        RECT 570.030 482.955 570.310 483.325 ;
        RECT 2008.450 162.675 2008.730 163.045 ;
        RECT 2008.520 82.870 2008.660 162.675 ;
        RECT 2008.520 82.730 2009.120 82.870 ;
        RECT 2008.980 2.400 2009.120 82.730 ;
        RECT 2008.770 -4.800 2009.330 2.400 ;
      LAYER via2 ;
        RECT 570.030 483.000 570.310 483.280 ;
        RECT 2008.450 162.720 2008.730 163.000 ;
      LAYER met3 ;
        RECT 568.830 483.290 569.210 483.300 ;
        RECT 570.005 483.290 570.335 483.305 ;
        RECT 568.830 482.990 570.335 483.290 ;
        RECT 568.830 482.980 569.210 482.990 ;
        RECT 570.005 482.975 570.335 482.990 ;
        RECT 568.830 163.010 569.210 163.020 ;
        RECT 2008.425 163.010 2008.755 163.025 ;
        RECT 568.830 162.710 2008.755 163.010 ;
        RECT 568.830 162.700 569.210 162.710 ;
        RECT 2008.425 162.695 2008.755 162.710 ;
      LAYER via3 ;
        RECT 568.860 482.980 569.180 483.300 ;
        RECT 568.860 162.700 569.180 163.020 ;
      LAYER met4 ;
        RECT 568.855 482.975 569.185 483.305 ;
        RECT 568.870 163.025 569.170 482.975 ;
        RECT 568.855 162.695 569.185 163.025 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.650 157.320 470.970 157.380 ;
        RECT 814.270 157.320 814.590 157.380 ;
        RECT 470.650 157.180 814.590 157.320 ;
        RECT 470.650 157.120 470.970 157.180 ;
        RECT 814.270 157.120 814.590 157.180 ;
      LAYER via ;
        RECT 470.680 157.120 470.940 157.380 ;
        RECT 814.300 157.120 814.560 157.380 ;
      LAYER met2 ;
        RECT 470.930 500.000 471.210 504.000 ;
        RECT 470.970 498.340 471.110 500.000 ;
        RECT 470.740 498.200 471.110 498.340 ;
        RECT 470.740 157.410 470.880 498.200 ;
        RECT 470.680 157.090 470.940 157.410 ;
        RECT 814.300 157.090 814.560 157.410 ;
        RECT 814.360 82.870 814.500 157.090 ;
        RECT 814.360 82.730 816.800 82.870 ;
        RECT 816.660 2.400 816.800 82.730 ;
        RECT 816.450 -4.800 817.010 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.670 500.000 571.950 504.000 ;
        RECT 571.710 498.965 571.850 500.000 ;
        RECT 571.640 498.595 571.920 498.965 ;
        RECT 2025.470 79.715 2025.750 80.085 ;
        RECT 2025.540 2.400 2025.680 79.715 ;
        RECT 2025.330 -4.800 2025.890 2.400 ;
      LAYER via2 ;
        RECT 571.640 498.640 571.920 498.920 ;
        RECT 2025.470 79.760 2025.750 80.040 ;
      LAYER met3 ;
        RECT 570.670 498.930 571.050 498.940 ;
        RECT 571.615 498.930 571.945 498.945 ;
        RECT 570.670 498.630 571.945 498.930 ;
        RECT 570.670 498.620 571.050 498.630 ;
        RECT 571.615 498.615 571.945 498.630 ;
        RECT 570.670 80.050 571.050 80.060 ;
        RECT 2025.445 80.050 2025.775 80.065 ;
        RECT 570.670 79.750 2025.775 80.050 ;
        RECT 570.670 79.740 571.050 79.750 ;
        RECT 2025.445 79.735 2025.775 79.750 ;
      LAYER via3 ;
        RECT 570.700 498.620 571.020 498.940 ;
        RECT 570.700 79.740 571.020 80.060 ;
      LAYER met4 ;
        RECT 570.695 498.615 571.025 498.945 ;
        RECT 570.710 80.065 571.010 498.615 ;
        RECT 570.695 79.735 571.025 80.065 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 472.160 573.090 472.220 ;
        RECT 575.530 472.160 575.850 472.220 ;
        RECT 572.770 472.020 575.850 472.160 ;
        RECT 572.770 471.960 573.090 472.020 ;
        RECT 575.530 471.960 575.850 472.020 ;
        RECT 575.530 170.920 575.850 170.980 ;
        RECT 2036.030 170.920 2036.350 170.980 ;
        RECT 575.530 170.780 2036.350 170.920 ;
        RECT 575.530 170.720 575.850 170.780 ;
        RECT 2036.030 170.720 2036.350 170.780 ;
        RECT 2036.030 20.300 2036.350 20.360 ;
        RECT 2042.010 20.300 2042.330 20.360 ;
        RECT 2036.030 20.160 2042.330 20.300 ;
        RECT 2036.030 20.100 2036.350 20.160 ;
        RECT 2042.010 20.100 2042.330 20.160 ;
      LAYER via ;
        RECT 572.800 471.960 573.060 472.220 ;
        RECT 575.560 471.960 575.820 472.220 ;
        RECT 575.560 170.720 575.820 170.980 ;
        RECT 2036.060 170.720 2036.320 170.980 ;
        RECT 2036.060 20.100 2036.320 20.360 ;
        RECT 2042.040 20.100 2042.300 20.360 ;
      LAYER met2 ;
        RECT 573.050 500.000 573.330 504.000 ;
        RECT 573.090 498.850 573.230 500.000 ;
        RECT 572.860 498.710 573.230 498.850 ;
        RECT 572.860 472.250 573.000 498.710 ;
        RECT 572.800 471.930 573.060 472.250 ;
        RECT 575.560 471.930 575.820 472.250 ;
        RECT 575.620 171.010 575.760 471.930 ;
        RECT 575.560 170.690 575.820 171.010 ;
        RECT 2036.060 170.690 2036.320 171.010 ;
        RECT 2036.120 20.390 2036.260 170.690 ;
        RECT 2036.060 20.070 2036.320 20.390 ;
        RECT 2042.040 20.070 2042.300 20.390 ;
        RECT 2042.100 2.400 2042.240 20.070 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.470 499.900 576.450 500.040 ;
        RECT 574.470 499.760 574.610 499.900 ;
        RECT 574.380 499.500 574.700 499.760 ;
        RECT 575.070 498.000 575.390 498.060 ;
        RECT 576.310 498.000 576.450 499.900 ;
        RECT 575.070 497.860 576.450 498.000 ;
        RECT 575.070 497.800 575.390 497.860 ;
        RECT 575.070 170.580 575.390 170.640 ;
        RECT 2056.270 170.580 2056.590 170.640 ;
        RECT 575.070 170.440 2056.590 170.580 ;
        RECT 575.070 170.380 575.390 170.440 ;
        RECT 2056.270 170.380 2056.590 170.440 ;
      LAYER via ;
        RECT 574.410 499.500 574.670 499.760 ;
        RECT 575.100 497.800 575.360 498.060 ;
        RECT 575.100 170.380 575.360 170.640 ;
        RECT 2056.300 170.380 2056.560 170.640 ;
      LAYER met2 ;
        RECT 574.430 500.000 574.710 504.000 ;
        RECT 574.470 499.790 574.610 500.000 ;
        RECT 574.410 499.470 574.670 499.790 ;
        RECT 575.100 497.770 575.360 498.090 ;
        RECT 575.160 170.670 575.300 497.770 ;
        RECT 575.100 170.350 575.360 170.670 ;
        RECT 2056.300 170.350 2056.560 170.670 ;
        RECT 2056.360 82.870 2056.500 170.350 ;
        RECT 2056.360 82.730 2058.800 82.870 ;
        RECT 2058.660 2.400 2058.800 82.730 ;
        RECT 2058.450 -4.800 2059.010 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 575.760 499.500 576.080 499.760 ;
        RECT 575.850 498.400 575.990 499.500 ;
        RECT 575.530 498.200 575.990 498.400 ;
        RECT 575.530 498.140 575.850 498.200 ;
        RECT 574.610 479.980 574.930 480.040 ;
        RECT 575.530 479.980 575.850 480.040 ;
        RECT 574.610 479.840 575.850 479.980 ;
        RECT 574.610 479.780 574.930 479.840 ;
        RECT 575.530 479.780 575.850 479.840 ;
        RECT 574.610 170.240 574.930 170.300 ;
        RECT 2070.070 170.240 2070.390 170.300 ;
        RECT 574.610 170.100 2070.390 170.240 ;
        RECT 574.610 170.040 574.930 170.100 ;
        RECT 2070.070 170.040 2070.390 170.100 ;
      LAYER via ;
        RECT 575.790 499.500 576.050 499.760 ;
        RECT 575.560 498.140 575.820 498.400 ;
        RECT 574.640 479.780 574.900 480.040 ;
        RECT 575.560 479.780 575.820 480.040 ;
        RECT 574.640 170.040 574.900 170.300 ;
        RECT 2070.100 170.040 2070.360 170.300 ;
      LAYER met2 ;
        RECT 575.810 500.000 576.090 504.000 ;
        RECT 575.850 499.790 575.990 500.000 ;
        RECT 575.790 499.470 576.050 499.790 ;
        RECT 575.560 498.110 575.820 498.430 ;
        RECT 575.620 480.070 575.760 498.110 ;
        RECT 574.640 479.750 574.900 480.070 ;
        RECT 575.560 479.750 575.820 480.070 ;
        RECT 574.700 170.330 574.840 479.750 ;
        RECT 574.640 170.010 574.900 170.330 ;
        RECT 2070.100 170.010 2070.360 170.330 ;
        RECT 2070.160 82.870 2070.300 170.010 ;
        RECT 2070.160 82.730 2075.360 82.870 ;
        RECT 2075.220 2.400 2075.360 82.730 ;
        RECT 2075.010 -4.800 2075.570 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 577.140 499.500 577.460 499.760 ;
        RECT 577.230 498.400 577.370 499.500 ;
        RECT 577.230 498.200 577.690 498.400 ;
        RECT 577.370 498.140 577.690 498.200 ;
        RECT 572.770 450.060 573.090 450.120 ;
        RECT 578.290 450.060 578.610 450.120 ;
        RECT 572.770 449.920 578.610 450.060 ;
        RECT 572.770 449.860 573.090 449.920 ;
        RECT 578.290 449.860 578.610 449.920 ;
        RECT 572.770 80.480 573.090 80.540 ;
        RECT 2091.690 80.480 2092.010 80.540 ;
        RECT 572.770 80.340 2092.010 80.480 ;
        RECT 572.770 80.280 573.090 80.340 ;
        RECT 2091.690 80.280 2092.010 80.340 ;
      LAYER via ;
        RECT 577.170 499.500 577.430 499.760 ;
        RECT 577.400 498.140 577.660 498.400 ;
        RECT 572.800 449.860 573.060 450.120 ;
        RECT 578.320 449.860 578.580 450.120 ;
        RECT 572.800 80.280 573.060 80.540 ;
        RECT 2091.720 80.280 2091.980 80.540 ;
      LAYER met2 ;
        RECT 577.190 500.000 577.470 504.000 ;
        RECT 577.230 499.790 577.370 500.000 ;
        RECT 577.170 499.470 577.430 499.790 ;
        RECT 577.400 498.110 577.660 498.430 ;
        RECT 577.460 477.090 577.600 498.110 ;
        RECT 577.460 476.950 578.520 477.090 ;
        RECT 578.380 450.150 578.520 476.950 ;
        RECT 572.800 449.830 573.060 450.150 ;
        RECT 578.320 449.830 578.580 450.150 ;
        RECT 572.860 80.570 573.000 449.830 ;
        RECT 572.800 80.250 573.060 80.570 ;
        RECT 2091.720 80.250 2091.980 80.570 ;
        RECT 2091.780 2.400 2091.920 80.250 ;
        RECT 2091.570 -4.800 2092.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 578.520 498.820 578.840 499.080 ;
        RECT 578.610 497.720 578.750 498.820 ;
        RECT 578.290 497.520 578.750 497.720 ;
        RECT 578.290 497.460 578.610 497.520 ;
      LAYER via ;
        RECT 578.550 498.820 578.810 499.080 ;
        RECT 578.320 497.460 578.580 497.720 ;
      LAYER met2 ;
        RECT 578.570 500.000 578.850 504.000 ;
        RECT 578.610 499.110 578.750 500.000 ;
        RECT 578.550 498.790 578.810 499.110 ;
        RECT 578.320 497.430 578.580 497.750 ;
        RECT 578.380 484.005 578.520 497.430 ;
        RECT 578.310 483.635 578.590 484.005 ;
        RECT 2104.590 453.715 2104.870 454.085 ;
        RECT 2104.660 82.870 2104.800 453.715 ;
        RECT 2104.660 82.730 2108.480 82.870 ;
        RECT 2108.340 2.400 2108.480 82.730 ;
        RECT 2108.130 -4.800 2108.690 2.400 ;
      LAYER via2 ;
        RECT 578.310 483.680 578.590 483.960 ;
        RECT 2104.590 453.760 2104.870 454.040 ;
      LAYER met3 ;
        RECT 578.285 483.980 578.615 483.985 ;
        RECT 578.030 483.970 578.615 483.980 ;
        RECT 578.030 483.670 578.840 483.970 ;
        RECT 578.030 483.660 578.615 483.670 ;
        RECT 578.285 483.655 578.615 483.660 ;
        RECT 578.030 454.050 578.410 454.060 ;
        RECT 2104.565 454.050 2104.895 454.065 ;
        RECT 578.030 453.750 2104.895 454.050 ;
        RECT 578.030 453.740 578.410 453.750 ;
        RECT 2104.565 453.735 2104.895 453.750 ;
      LAYER via3 ;
        RECT 578.060 483.660 578.380 483.980 ;
        RECT 578.060 453.740 578.380 454.060 ;
      LAYER met4 ;
        RECT 578.055 483.655 578.385 483.985 ;
        RECT 578.070 454.065 578.370 483.655 ;
        RECT 578.055 453.735 578.385 454.065 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.900 499.500 580.220 499.760 ;
        RECT 579.990 498.340 580.130 499.500 ;
        RECT 579.990 498.200 580.820 498.340 ;
        RECT 579.670 497.660 579.990 497.720 ;
        RECT 580.680 497.660 580.820 498.200 ;
        RECT 579.670 497.520 580.820 497.660 ;
        RECT 579.670 497.460 579.990 497.520 ;
        RECT 579.670 80.140 579.990 80.200 ;
        RECT 2118.830 80.140 2119.150 80.200 ;
        RECT 579.670 80.000 2119.150 80.140 ;
        RECT 579.670 79.940 579.990 80.000 ;
        RECT 2118.830 79.940 2119.150 80.000 ;
        RECT 2118.830 19.280 2119.150 19.340 ;
        RECT 2124.810 19.280 2125.130 19.340 ;
        RECT 2118.830 19.140 2125.130 19.280 ;
        RECT 2118.830 19.080 2119.150 19.140 ;
        RECT 2124.810 19.080 2125.130 19.140 ;
      LAYER via ;
        RECT 579.930 499.500 580.190 499.760 ;
        RECT 579.700 497.460 579.960 497.720 ;
        RECT 579.700 79.940 579.960 80.200 ;
        RECT 2118.860 79.940 2119.120 80.200 ;
        RECT 2118.860 19.080 2119.120 19.340 ;
        RECT 2124.840 19.080 2125.100 19.340 ;
      LAYER met2 ;
        RECT 579.950 500.000 580.230 504.000 ;
        RECT 579.990 499.790 580.130 500.000 ;
        RECT 579.930 499.470 580.190 499.790 ;
        RECT 579.700 497.430 579.960 497.750 ;
        RECT 579.760 80.230 579.900 497.430 ;
        RECT 579.700 79.910 579.960 80.230 ;
        RECT 2118.860 79.910 2119.120 80.230 ;
        RECT 2118.920 19.370 2119.060 79.910 ;
        RECT 2118.860 19.050 2119.120 19.370 ;
        RECT 2124.840 19.050 2125.100 19.370 ;
        RECT 2124.900 2.400 2125.040 19.050 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.280 499.160 581.600 499.420 ;
        RECT 581.370 498.400 581.510 499.160 ;
        RECT 581.370 498.200 581.830 498.400 ;
        RECT 581.510 498.140 581.830 498.200 ;
        RECT 580.130 472.840 580.450 472.900 ;
        RECT 581.510 472.840 581.830 472.900 ;
        RECT 580.130 472.700 581.830 472.840 ;
        RECT 580.130 472.640 580.450 472.700 ;
        RECT 581.510 472.640 581.830 472.700 ;
        RECT 580.130 169.900 580.450 169.960 ;
        RECT 2139.070 169.900 2139.390 169.960 ;
        RECT 580.130 169.760 2139.390 169.900 ;
        RECT 580.130 169.700 580.450 169.760 ;
        RECT 2139.070 169.700 2139.390 169.760 ;
      LAYER via ;
        RECT 581.310 499.160 581.570 499.420 ;
        RECT 581.540 498.140 581.800 498.400 ;
        RECT 580.160 472.640 580.420 472.900 ;
        RECT 581.540 472.640 581.800 472.900 ;
        RECT 580.160 169.700 580.420 169.960 ;
        RECT 2139.100 169.700 2139.360 169.960 ;
      LAYER met2 ;
        RECT 581.330 500.000 581.610 504.000 ;
        RECT 581.370 499.450 581.510 500.000 ;
        RECT 581.310 499.130 581.570 499.450 ;
        RECT 581.540 498.110 581.800 498.430 ;
        RECT 581.600 472.930 581.740 498.110 ;
        RECT 580.160 472.610 580.420 472.930 ;
        RECT 581.540 472.610 581.800 472.930 ;
        RECT 580.220 169.990 580.360 472.610 ;
        RECT 580.160 169.670 580.420 169.990 ;
        RECT 2139.100 169.670 2139.360 169.990 ;
        RECT 2139.160 82.870 2139.300 169.670 ;
        RECT 2139.160 82.730 2141.600 82.870 ;
        RECT 2141.460 2.400 2141.600 82.730 ;
        RECT 2141.250 -4.800 2141.810 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 169.560 580.910 169.620 ;
        RECT 2152.870 169.560 2153.190 169.620 ;
        RECT 580.590 169.420 2153.190 169.560 ;
        RECT 580.590 169.360 580.910 169.420 ;
        RECT 2152.870 169.360 2153.190 169.420 ;
      LAYER via ;
        RECT 580.620 169.360 580.880 169.620 ;
        RECT 2152.900 169.360 2153.160 169.620 ;
      LAYER met2 ;
        RECT 582.710 500.000 582.990 504.000 ;
        RECT 582.750 499.645 582.890 500.000 ;
        RECT 582.680 499.275 582.960 499.645 ;
        RECT 580.610 497.235 580.890 497.605 ;
        RECT 580.680 169.650 580.820 497.235 ;
        RECT 580.620 169.330 580.880 169.650 ;
        RECT 2152.900 169.330 2153.160 169.650 ;
        RECT 2152.960 82.870 2153.100 169.330 ;
        RECT 2152.960 82.730 2158.160 82.870 ;
        RECT 2158.020 2.400 2158.160 82.730 ;
        RECT 2157.810 -4.800 2158.370 2.400 ;
      LAYER via2 ;
        RECT 582.680 499.320 582.960 499.600 ;
        RECT 580.610 497.280 580.890 497.560 ;
      LAYER met3 ;
        RECT 582.655 499.295 582.985 499.625 ;
        RECT 580.585 497.570 580.915 497.585 ;
        RECT 582.670 497.570 582.970 499.295 ;
        RECT 580.585 497.270 582.970 497.570 ;
        RECT 580.585 497.255 580.915 497.270 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.040 499.500 584.360 499.760 ;
        RECT 584.130 499.360 584.270 499.500 ;
        RECT 584.130 499.220 584.960 499.360 ;
        RECT 583.810 498.000 584.130 498.060 ;
        RECT 584.820 498.000 584.960 499.220 ;
        RECT 583.810 497.860 584.960 498.000 ;
        RECT 583.810 497.800 584.130 497.860 ;
      LAYER via ;
        RECT 584.070 499.500 584.330 499.760 ;
        RECT 583.840 497.800 584.100 498.060 ;
      LAYER met2 ;
        RECT 584.090 500.000 584.370 504.000 ;
        RECT 584.130 499.790 584.270 500.000 ;
        RECT 584.070 499.470 584.330 499.790 ;
        RECT 583.840 497.770 584.100 498.090 ;
        RECT 583.900 487.405 584.040 497.770 ;
        RECT 583.830 487.035 584.110 487.405 ;
        RECT 2174.050 178.315 2174.330 178.685 ;
        RECT 2174.120 82.870 2174.260 178.315 ;
        RECT 2174.120 82.730 2174.720 82.870 ;
        RECT 2174.580 2.400 2174.720 82.730 ;
        RECT 2174.370 -4.800 2174.930 2.400 ;
      LAYER via2 ;
        RECT 583.830 487.080 584.110 487.360 ;
        RECT 2174.050 178.360 2174.330 178.640 ;
      LAYER met3 ;
        RECT 583.805 487.370 584.135 487.385 ;
        RECT 584.470 487.370 584.850 487.380 ;
        RECT 583.805 487.070 584.850 487.370 ;
        RECT 583.805 487.055 584.135 487.070 ;
        RECT 584.470 487.060 584.850 487.070 ;
        RECT 584.470 178.650 584.850 178.660 ;
        RECT 2174.025 178.650 2174.355 178.665 ;
        RECT 584.470 178.350 2174.355 178.650 ;
        RECT 584.470 178.340 584.850 178.350 ;
        RECT 2174.025 178.335 2174.355 178.350 ;
      LAYER via3 ;
        RECT 584.500 487.060 584.820 487.380 ;
        RECT 584.500 178.340 584.820 178.660 ;
      LAYER met4 ;
        RECT 584.495 487.055 584.825 487.385 ;
        RECT 584.510 178.665 584.810 487.055 ;
        RECT 584.495 178.335 584.825 178.665 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 471.110 472.840 471.430 472.900 ;
        RECT 472.030 472.840 472.350 472.900 ;
        RECT 471.110 472.700 472.350 472.840 ;
        RECT 471.110 472.640 471.430 472.700 ;
        RECT 472.030 472.640 472.350 472.700 ;
        RECT 471.110 205.940 471.430 206.000 ;
        RECT 828.070 205.940 828.390 206.000 ;
        RECT 471.110 205.800 828.390 205.940 ;
        RECT 471.110 205.740 471.430 205.800 ;
        RECT 828.070 205.740 828.390 205.800 ;
      LAYER via ;
        RECT 471.140 472.640 471.400 472.900 ;
        RECT 472.060 472.640 472.320 472.900 ;
        RECT 471.140 205.740 471.400 206.000 ;
        RECT 828.100 205.740 828.360 206.000 ;
      LAYER met2 ;
        RECT 472.310 500.000 472.590 504.000 ;
        RECT 472.350 499.020 472.490 500.000 ;
        RECT 472.120 498.880 472.490 499.020 ;
        RECT 472.120 472.930 472.260 498.880 ;
        RECT 471.140 472.610 471.400 472.930 ;
        RECT 472.060 472.610 472.320 472.930 ;
        RECT 471.200 206.030 471.340 472.610 ;
        RECT 471.140 205.710 471.400 206.030 ;
        RECT 828.100 205.710 828.360 206.030 ;
        RECT 828.160 82.870 828.300 205.710 ;
        RECT 828.160 82.730 833.360 82.870 ;
        RECT 833.220 2.400 833.360 82.730 ;
        RECT 833.010 -4.800 833.570 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.470 500.000 585.750 504.000 ;
        RECT 585.510 499.815 585.650 500.000 ;
        RECT 585.440 499.445 585.720 499.815 ;
        RECT 2187.390 177.635 2187.670 178.005 ;
        RECT 2187.460 82.870 2187.600 177.635 ;
        RECT 2187.460 82.730 2191.280 82.870 ;
        RECT 2191.140 2.400 2191.280 82.730 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
      LAYER via2 ;
        RECT 585.440 499.490 585.720 499.770 ;
        RECT 2187.390 177.680 2187.670 177.960 ;
      LAYER met3 ;
        RECT 585.415 499.620 585.745 499.795 ;
        RECT 585.390 499.610 585.770 499.620 ;
        RECT 585.390 499.310 586.030 499.610 ;
        RECT 585.390 499.300 585.770 499.310 ;
        RECT 585.390 177.970 585.770 177.980 ;
        RECT 2187.365 177.970 2187.695 177.985 ;
        RECT 585.390 177.670 2187.695 177.970 ;
        RECT 585.390 177.660 585.770 177.670 ;
        RECT 2187.365 177.655 2187.695 177.670 ;
      LAYER via3 ;
        RECT 585.420 499.300 585.740 499.620 ;
        RECT 585.420 177.660 585.740 177.980 ;
      LAYER met4 ;
        RECT 585.415 499.295 585.745 499.625 ;
        RECT 585.430 177.985 585.730 499.295 ;
        RECT 585.415 177.655 585.745 177.985 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.800 499.500 587.120 499.760 ;
        RECT 586.890 498.060 587.030 499.500 ;
        RECT 586.890 497.860 587.350 498.060 ;
        RECT 587.030 497.800 587.350 497.860 ;
        RECT 587.490 177.040 587.810 177.100 ;
        RECT 2201.630 177.040 2201.950 177.100 ;
        RECT 587.490 176.900 2201.950 177.040 ;
        RECT 587.490 176.840 587.810 176.900 ;
        RECT 2201.630 176.840 2201.950 176.900 ;
        RECT 2201.630 19.280 2201.950 19.340 ;
        RECT 2207.610 19.280 2207.930 19.340 ;
        RECT 2201.630 19.140 2207.930 19.280 ;
        RECT 2201.630 19.080 2201.950 19.140 ;
        RECT 2207.610 19.080 2207.930 19.140 ;
      LAYER via ;
        RECT 586.830 499.500 587.090 499.760 ;
        RECT 587.060 497.800 587.320 498.060 ;
        RECT 587.520 176.840 587.780 177.100 ;
        RECT 2201.660 176.840 2201.920 177.100 ;
        RECT 2201.660 19.080 2201.920 19.340 ;
        RECT 2207.640 19.080 2207.900 19.340 ;
      LAYER met2 ;
        RECT 586.850 500.000 587.130 504.000 ;
        RECT 586.890 499.790 587.030 500.000 ;
        RECT 586.830 499.470 587.090 499.790 ;
        RECT 587.060 497.770 587.320 498.090 ;
        RECT 587.120 473.010 587.260 497.770 ;
        RECT 587.120 472.870 587.720 473.010 ;
        RECT 587.580 177.130 587.720 472.870 ;
        RECT 587.520 176.810 587.780 177.130 ;
        RECT 2201.660 176.810 2201.920 177.130 ;
        RECT 2201.720 19.370 2201.860 176.810 ;
        RECT 2201.660 19.050 2201.920 19.370 ;
        RECT 2207.640 19.050 2207.900 19.370 ;
        RECT 2207.700 2.400 2207.840 19.050 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.180 500.520 588.500 500.780 ;
        RECT 588.270 499.020 588.410 500.520 ;
        RECT 588.040 498.880 588.410 499.020 ;
        RECT 586.570 497.320 586.890 497.380 ;
        RECT 588.040 497.320 588.180 498.880 ;
        RECT 586.570 497.180 588.180 497.320 ;
        RECT 586.570 497.120 586.890 497.180 ;
        RECT 587.030 176.700 587.350 176.760 ;
        RECT 2221.870 176.700 2222.190 176.760 ;
        RECT 587.030 176.560 2222.190 176.700 ;
        RECT 587.030 176.500 587.350 176.560 ;
        RECT 2221.870 176.500 2222.190 176.560 ;
      LAYER via ;
        RECT 588.210 500.520 588.470 500.780 ;
        RECT 586.600 497.120 586.860 497.380 ;
        RECT 587.060 176.500 587.320 176.760 ;
        RECT 2221.900 176.500 2222.160 176.760 ;
      LAYER met2 ;
        RECT 588.230 500.810 588.510 504.000 ;
        RECT 588.210 500.490 588.510 500.810 ;
        RECT 588.230 500.000 588.510 500.490 ;
        RECT 586.600 497.090 586.860 497.410 ;
        RECT 586.660 472.330 586.800 497.090 ;
        RECT 586.660 472.190 587.260 472.330 ;
        RECT 587.120 176.790 587.260 472.190 ;
        RECT 587.060 176.470 587.320 176.790 ;
        RECT 2221.900 176.470 2222.160 176.790 ;
        RECT 2221.960 82.870 2222.100 176.470 ;
        RECT 2221.960 82.730 2224.400 82.870 ;
        RECT 2224.260 2.400 2224.400 82.730 ;
        RECT 2224.050 -4.800 2224.610 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 589.560 499.500 589.880 499.760 ;
        RECT 589.650 498.400 589.790 499.500 ;
        RECT 589.330 498.200 589.790 498.400 ;
        RECT 589.330 498.140 589.650 498.200 ;
        RECT 586.570 471.820 586.890 471.880 ;
        RECT 589.330 471.820 589.650 471.880 ;
        RECT 586.570 471.680 589.650 471.820 ;
        RECT 586.570 471.620 586.890 471.680 ;
        RECT 589.330 471.620 589.650 471.680 ;
        RECT 586.570 169.220 586.890 169.280 ;
        RECT 2235.670 169.220 2235.990 169.280 ;
        RECT 586.570 169.080 2235.990 169.220 ;
        RECT 586.570 169.020 586.890 169.080 ;
        RECT 2235.670 169.020 2235.990 169.080 ;
      LAYER via ;
        RECT 589.590 499.500 589.850 499.760 ;
        RECT 589.360 498.140 589.620 498.400 ;
        RECT 586.600 471.620 586.860 471.880 ;
        RECT 589.360 471.620 589.620 471.880 ;
        RECT 586.600 169.020 586.860 169.280 ;
        RECT 2235.700 169.020 2235.960 169.280 ;
      LAYER met2 ;
        RECT 589.610 500.000 589.890 504.000 ;
        RECT 589.650 499.790 589.790 500.000 ;
        RECT 589.590 499.470 589.850 499.790 ;
        RECT 589.360 498.110 589.620 498.430 ;
        RECT 589.420 471.910 589.560 498.110 ;
        RECT 586.600 471.590 586.860 471.910 ;
        RECT 589.360 471.590 589.620 471.910 ;
        RECT 586.660 169.310 586.800 471.590 ;
        RECT 586.600 168.990 586.860 169.310 ;
        RECT 2235.700 168.990 2235.960 169.310 ;
        RECT 2235.760 82.870 2235.900 168.990 ;
        RECT 2235.760 82.730 2240.960 82.870 ;
        RECT 2240.820 2.400 2240.960 82.730 ;
        RECT 2240.610 -4.800 2241.170 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.940 499.160 591.260 499.420 ;
        RECT 591.030 498.740 591.170 499.160 ;
        RECT 591.030 498.540 591.490 498.740 ;
        RECT 591.170 498.480 591.490 498.540 ;
      LAYER via ;
        RECT 590.970 499.160 591.230 499.420 ;
        RECT 591.200 498.480 591.460 498.740 ;
      LAYER met2 ;
        RECT 590.990 500.000 591.270 504.000 ;
        RECT 591.030 499.450 591.170 500.000 ;
        RECT 590.970 499.130 591.230 499.450 ;
        RECT 591.190 498.595 591.470 498.965 ;
        RECT 591.200 498.450 591.460 498.595 ;
        RECT 2256.850 176.955 2257.130 177.325 ;
        RECT 2256.920 82.870 2257.060 176.955 ;
        RECT 2256.920 82.730 2257.520 82.870 ;
        RECT 2257.380 2.400 2257.520 82.730 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
      LAYER via2 ;
        RECT 591.190 498.640 591.470 498.920 ;
        RECT 2256.850 177.000 2257.130 177.280 ;
      LAYER met3 ;
        RECT 591.165 498.940 591.495 498.945 ;
        RECT 590.910 498.930 591.495 498.940 ;
        RECT 590.710 498.630 591.495 498.930 ;
        RECT 590.910 498.620 591.495 498.630 ;
        RECT 591.165 498.615 591.495 498.620 ;
        RECT 590.910 177.290 591.290 177.300 ;
        RECT 2256.825 177.290 2257.155 177.305 ;
        RECT 590.910 176.990 2257.155 177.290 ;
        RECT 590.910 176.980 591.290 176.990 ;
        RECT 2256.825 176.975 2257.155 176.990 ;
      LAYER via3 ;
        RECT 590.940 498.620 591.260 498.940 ;
        RECT 590.940 176.980 591.260 177.300 ;
      LAYER met4 ;
        RECT 590.935 498.615 591.265 498.945 ;
        RECT 590.950 177.305 591.250 498.615 ;
        RECT 590.935 176.975 591.265 177.305 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.370 500.000 592.650 504.000 ;
        RECT 592.410 499.815 592.550 500.000 ;
        RECT 592.340 499.445 592.620 499.815 ;
        RECT 2270.190 176.275 2270.470 176.645 ;
        RECT 2270.260 82.870 2270.400 176.275 ;
        RECT 2270.260 82.730 2274.080 82.870 ;
        RECT 2273.940 2.400 2274.080 82.730 ;
        RECT 2273.730 -4.800 2274.290 2.400 ;
      LAYER via2 ;
        RECT 592.340 499.490 592.620 499.770 ;
        RECT 2270.190 176.320 2270.470 176.600 ;
      LAYER met3 ;
        RECT 592.315 499.465 592.645 499.795 ;
        RECT 589.990 498.250 590.370 498.260 ;
        RECT 592.330 498.250 592.630 499.465 ;
        RECT 589.990 497.950 592.630 498.250 ;
        RECT 589.990 497.940 590.370 497.950 ;
        RECT 589.990 176.610 590.370 176.620 ;
        RECT 2270.165 176.610 2270.495 176.625 ;
        RECT 589.990 176.310 2270.495 176.610 ;
        RECT 589.990 176.300 590.370 176.310 ;
        RECT 2270.165 176.295 2270.495 176.310 ;
      LAYER via3 ;
        RECT 590.020 497.940 590.340 498.260 ;
        RECT 590.020 176.300 590.340 176.620 ;
      LAYER met4 ;
        RECT 590.015 497.935 590.345 498.265 ;
        RECT 590.030 176.625 590.330 497.935 ;
        RECT 590.015 176.295 590.345 176.625 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.700 499.160 594.020 499.420 ;
        RECT 593.790 497.720 593.930 499.160 ;
        RECT 593.790 497.520 594.250 497.720 ;
        RECT 593.930 497.460 594.250 497.520 ;
        RECT 593.930 484.740 594.250 484.800 ;
        RECT 595.770 484.740 596.090 484.800 ;
        RECT 593.930 484.600 596.090 484.740 ;
        RECT 593.930 484.540 594.250 484.600 ;
        RECT 595.770 484.540 596.090 484.600 ;
        RECT 595.770 204.240 596.090 204.300 ;
        RECT 2284.430 204.240 2284.750 204.300 ;
        RECT 595.770 204.100 2284.750 204.240 ;
        RECT 595.770 204.040 596.090 204.100 ;
        RECT 2284.430 204.040 2284.750 204.100 ;
        RECT 2284.430 18.600 2284.750 18.660 ;
        RECT 2290.410 18.600 2290.730 18.660 ;
        RECT 2284.430 18.460 2290.730 18.600 ;
        RECT 2284.430 18.400 2284.750 18.460 ;
        RECT 2290.410 18.400 2290.730 18.460 ;
      LAYER via ;
        RECT 593.730 499.160 593.990 499.420 ;
        RECT 593.960 497.460 594.220 497.720 ;
        RECT 593.960 484.540 594.220 484.800 ;
        RECT 595.800 484.540 596.060 484.800 ;
        RECT 595.800 204.040 596.060 204.300 ;
        RECT 2284.460 204.040 2284.720 204.300 ;
        RECT 2284.460 18.400 2284.720 18.660 ;
        RECT 2290.440 18.400 2290.700 18.660 ;
      LAYER met2 ;
        RECT 593.750 500.000 594.030 504.000 ;
        RECT 593.790 499.450 593.930 500.000 ;
        RECT 593.730 499.130 593.990 499.450 ;
        RECT 593.960 497.430 594.220 497.750 ;
        RECT 594.020 484.830 594.160 497.430 ;
        RECT 593.960 484.510 594.220 484.830 ;
        RECT 595.800 484.510 596.060 484.830 ;
        RECT 595.860 204.330 596.000 484.510 ;
        RECT 595.800 204.010 596.060 204.330 ;
        RECT 2284.460 204.010 2284.720 204.330 ;
        RECT 2284.520 18.690 2284.660 204.010 ;
        RECT 2284.460 18.370 2284.720 18.690 ;
        RECT 2290.440 18.370 2290.700 18.690 ;
        RECT 2290.500 2.400 2290.640 18.370 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 595.310 203.900 595.630 203.960 ;
        RECT 2304.670 203.900 2304.990 203.960 ;
        RECT 595.310 203.760 2304.990 203.900 ;
        RECT 595.310 203.700 595.630 203.760 ;
        RECT 2304.670 203.700 2304.990 203.760 ;
      LAYER via ;
        RECT 595.340 203.700 595.600 203.960 ;
        RECT 2304.700 203.700 2304.960 203.960 ;
      LAYER met2 ;
        RECT 595.130 500.000 595.410 504.000 ;
        RECT 595.170 498.680 595.310 500.000 ;
        RECT 595.170 498.540 595.540 498.680 ;
        RECT 595.400 203.990 595.540 498.540 ;
        RECT 595.340 203.670 595.600 203.990 ;
        RECT 2304.700 203.670 2304.960 203.990 ;
        RECT 2304.760 82.870 2304.900 203.670 ;
        RECT 2304.760 82.730 2307.200 82.870 ;
        RECT 2307.060 2.400 2307.200 82.730 ;
        RECT 2306.850 -4.800 2307.410 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.460 498.820 596.780 499.080 ;
        RECT 596.550 498.680 596.690 498.820 ;
        RECT 596.550 498.540 598.300 498.680 ;
        RECT 598.160 498.400 598.300 498.540 ;
        RECT 598.070 498.140 598.390 498.400 ;
        RECT 594.850 486.440 595.170 486.500 ;
        RECT 598.070 486.440 598.390 486.500 ;
        RECT 594.850 486.300 598.390 486.440 ;
        RECT 594.850 486.240 595.170 486.300 ;
        RECT 598.070 486.240 598.390 486.300 ;
        RECT 594.850 120.600 595.170 120.660 ;
        RECT 2318.470 120.600 2318.790 120.660 ;
        RECT 594.850 120.460 2318.790 120.600 ;
        RECT 594.850 120.400 595.170 120.460 ;
        RECT 2318.470 120.400 2318.790 120.460 ;
      LAYER via ;
        RECT 596.490 498.820 596.750 499.080 ;
        RECT 598.100 498.140 598.360 498.400 ;
        RECT 594.880 486.240 595.140 486.500 ;
        RECT 598.100 486.240 598.360 486.500 ;
        RECT 594.880 120.400 595.140 120.660 ;
        RECT 2318.500 120.400 2318.760 120.660 ;
      LAYER met2 ;
        RECT 596.510 500.000 596.790 504.000 ;
        RECT 596.550 499.110 596.690 500.000 ;
        RECT 596.490 498.790 596.750 499.110 ;
        RECT 598.100 498.110 598.360 498.430 ;
        RECT 598.160 486.530 598.300 498.110 ;
        RECT 594.880 486.210 595.140 486.530 ;
        RECT 598.100 486.210 598.360 486.530 ;
        RECT 594.940 120.690 595.080 486.210 ;
        RECT 594.880 120.370 595.140 120.690 ;
        RECT 2318.500 120.370 2318.760 120.690 ;
        RECT 2318.560 82.870 2318.700 120.370 ;
        RECT 2318.560 82.730 2323.760 82.870 ;
        RECT 2323.620 2.400 2323.760 82.730 ;
        RECT 2323.410 -4.800 2323.970 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 597.840 499.500 598.160 499.760 ;
        RECT 597.930 499.360 598.070 499.500 ;
        RECT 597.930 499.220 598.300 499.360 ;
        RECT 598.160 499.080 598.300 499.220 ;
        RECT 598.070 498.820 598.390 499.080 ;
      LAYER via ;
        RECT 597.870 499.500 598.130 499.760 ;
        RECT 598.100 498.820 598.360 499.080 ;
      LAYER met2 ;
        RECT 597.890 500.000 598.170 504.000 ;
        RECT 597.930 499.790 598.070 500.000 ;
        RECT 597.870 499.470 598.130 499.790 ;
        RECT 598.100 498.965 598.360 499.110 ;
        RECT 598.090 498.595 598.370 498.965 ;
        RECT 2339.650 161.995 2339.930 162.365 ;
        RECT 2339.720 82.870 2339.860 161.995 ;
        RECT 2339.720 82.730 2340.320 82.870 ;
        RECT 2340.180 2.400 2340.320 82.730 ;
        RECT 2339.970 -4.800 2340.530 2.400 ;
      LAYER via2 ;
        RECT 598.090 498.640 598.370 498.920 ;
        RECT 2339.650 162.040 2339.930 162.320 ;
      LAYER met3 ;
        RECT 598.065 498.940 598.395 498.945 ;
        RECT 598.065 498.930 598.650 498.940 ;
        RECT 598.065 498.630 598.850 498.930 ;
        RECT 598.065 498.620 598.650 498.630 ;
        RECT 598.065 498.615 598.395 498.620 ;
        RECT 598.270 162.330 598.650 162.340 ;
        RECT 2339.625 162.330 2339.955 162.345 ;
        RECT 598.270 162.030 2339.955 162.330 ;
        RECT 598.270 162.020 598.650 162.030 ;
        RECT 2339.625 162.015 2339.955 162.030 ;
      LAYER via3 ;
        RECT 598.300 498.620 598.620 498.940 ;
        RECT 598.300 162.020 598.620 162.340 ;
      LAYER met4 ;
        RECT 598.295 498.615 598.625 498.945 ;
        RECT 598.310 162.345 598.610 498.615 ;
        RECT 598.295 162.015 598.625 162.345 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 473.640 499.500 473.960 499.760 ;
        RECT 473.730 499.080 473.870 499.500 ;
        RECT 473.410 498.880 473.870 499.080 ;
        RECT 473.410 498.820 473.730 498.880 ;
      LAYER via ;
        RECT 473.670 499.500 473.930 499.760 ;
        RECT 473.440 498.820 473.700 499.080 ;
      LAYER met2 ;
        RECT 473.690 500.000 473.970 504.000 ;
        RECT 473.730 499.790 473.870 500.000 ;
        RECT 473.670 499.470 473.930 499.790 ;
        RECT 473.440 498.965 473.700 499.110 ;
        RECT 473.430 498.595 473.710 498.965 ;
        RECT 849.250 203.475 849.530 203.845 ;
        RECT 849.320 82.870 849.460 203.475 ;
        RECT 849.320 82.730 849.920 82.870 ;
        RECT 849.780 2.400 849.920 82.730 ;
        RECT 849.570 -4.800 850.130 2.400 ;
      LAYER via2 ;
        RECT 473.430 498.640 473.710 498.920 ;
        RECT 849.250 203.520 849.530 203.800 ;
      LAYER met3 ;
        RECT 473.405 498.940 473.735 498.945 ;
        RECT 473.150 498.930 473.735 498.940 ;
        RECT 472.950 498.630 473.735 498.930 ;
        RECT 473.150 498.620 473.735 498.630 ;
        RECT 473.405 498.615 473.735 498.620 ;
        RECT 473.150 203.810 473.530 203.820 ;
        RECT 849.225 203.810 849.555 203.825 ;
        RECT 473.150 203.510 849.555 203.810 ;
        RECT 473.150 203.500 473.530 203.510 ;
        RECT 849.225 203.495 849.555 203.510 ;
      LAYER via3 ;
        RECT 473.180 498.620 473.500 498.940 ;
        RECT 473.180 203.500 473.500 203.820 ;
      LAYER met4 ;
        RECT 473.175 498.615 473.505 498.945 ;
        RECT 473.190 203.825 473.490 498.615 ;
        RECT 473.175 203.495 473.505 203.825 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 461.680 499.500 462.000 499.760 ;
        RECT 461.770 498.400 461.910 499.500 ;
        RECT 461.450 498.200 461.910 498.400 ;
        RECT 461.450 498.140 461.770 498.200 ;
      LAYER via ;
        RECT 461.710 499.500 461.970 499.760 ;
        RECT 461.480 498.140 461.740 498.400 ;
      LAYER met2 ;
        RECT 461.730 500.000 462.010 504.000 ;
        RECT 461.770 499.790 461.910 500.000 ;
        RECT 461.710 499.470 461.970 499.790 ;
        RECT 461.480 498.170 461.740 498.430 ;
        RECT 461.080 498.110 461.740 498.170 ;
        RECT 461.080 498.030 461.680 498.110 ;
        RECT 461.080 490.805 461.220 498.030 ;
        RECT 461.010 490.435 461.290 490.805 ;
        RECT 703.890 204.155 704.170 204.525 ;
        RECT 703.960 82.870 704.100 204.155 ;
        RECT 703.960 82.730 706.400 82.870 ;
        RECT 706.260 2.400 706.400 82.730 ;
        RECT 706.050 -4.800 706.610 2.400 ;
      LAYER via2 ;
        RECT 461.010 490.480 461.290 490.760 ;
        RECT 703.890 204.200 704.170 204.480 ;
      LAYER met3 ;
        RECT 456.590 490.770 456.970 490.780 ;
        RECT 460.985 490.770 461.315 490.785 ;
        RECT 456.590 490.470 461.315 490.770 ;
        RECT 456.590 490.460 456.970 490.470 ;
        RECT 460.985 490.455 461.315 490.470 ;
        RECT 456.590 204.490 456.970 204.500 ;
        RECT 703.865 204.490 704.195 204.505 ;
        RECT 456.590 204.190 704.195 204.490 ;
        RECT 456.590 204.180 456.970 204.190 ;
        RECT 703.865 204.175 704.195 204.190 ;
      LAYER via3 ;
        RECT 456.620 490.460 456.940 490.780 ;
        RECT 456.620 204.180 456.940 204.500 ;
      LAYER met4 ;
        RECT 456.615 490.455 456.945 490.785 ;
        RECT 456.630 204.505 456.930 490.455 ;
        RECT 456.615 204.175 456.945 204.505 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 599.680 499.160 600.000 499.420 ;
        RECT 599.770 498.400 599.910 499.160 ;
        RECT 599.450 498.200 599.910 498.400 ;
        RECT 599.450 498.140 599.770 498.200 ;
      LAYER via ;
        RECT 599.710 499.160 599.970 499.420 ;
        RECT 599.480 498.140 599.740 498.400 ;
      LAYER met2 ;
        RECT 599.730 500.000 600.010 504.000 ;
        RECT 599.770 499.450 599.910 500.000 ;
        RECT 599.710 499.130 599.970 499.450 ;
        RECT 599.480 498.110 599.740 498.430 ;
        RECT 599.540 480.605 599.680 498.110 ;
        RECT 599.470 480.235 599.750 480.605 ;
        RECT 2359.890 480.235 2360.170 480.605 ;
        RECT 2359.960 82.870 2360.100 480.235 ;
        RECT 2359.960 82.730 2362.400 82.870 ;
        RECT 2362.260 2.400 2362.400 82.730 ;
        RECT 2362.050 -4.800 2362.610 2.400 ;
      LAYER via2 ;
        RECT 599.470 480.280 599.750 480.560 ;
        RECT 2359.890 480.280 2360.170 480.560 ;
      LAYER met3 ;
        RECT 599.445 480.570 599.775 480.585 ;
        RECT 2359.865 480.570 2360.195 480.585 ;
        RECT 599.445 480.270 2360.195 480.570 ;
        RECT 599.445 480.255 599.775 480.270 ;
        RECT 2359.865 480.255 2360.195 480.270 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 86.940 602.070 87.000 ;
        RECT 2373.670 86.940 2373.990 87.000 ;
        RECT 601.750 86.800 2373.990 86.940 ;
        RECT 601.750 86.740 602.070 86.800 ;
        RECT 2373.670 86.740 2373.990 86.800 ;
      LAYER via ;
        RECT 601.780 86.740 602.040 87.000 ;
        RECT 2373.700 86.740 2373.960 87.000 ;
      LAYER met2 ;
        RECT 601.110 500.000 601.390 504.000 ;
        RECT 601.150 498.680 601.290 500.000 ;
        RECT 601.150 498.540 601.520 498.680 ;
        RECT 601.380 469.270 601.520 498.540 ;
        RECT 601.380 469.130 601.980 469.270 ;
        RECT 601.840 87.030 601.980 469.130 ;
        RECT 601.780 86.710 602.040 87.030 ;
        RECT 2373.700 86.710 2373.960 87.030 ;
        RECT 2373.760 82.870 2373.900 86.710 ;
        RECT 2373.760 82.730 2378.960 82.870 ;
        RECT 2378.820 2.400 2378.960 82.730 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 602.440 499.500 602.760 499.760 ;
        RECT 602.530 498.740 602.670 499.500 ;
        RECT 602.530 498.540 602.990 498.740 ;
        RECT 602.670 498.480 602.990 498.540 ;
        RECT 602.670 148.140 602.990 148.200 ;
        RECT 2394.830 148.140 2395.150 148.200 ;
        RECT 602.670 148.000 2395.150 148.140 ;
        RECT 602.670 147.940 602.990 148.000 ;
        RECT 2394.830 147.940 2395.150 148.000 ;
      LAYER via ;
        RECT 602.470 499.500 602.730 499.760 ;
        RECT 602.700 498.480 602.960 498.740 ;
        RECT 602.700 147.940 602.960 148.200 ;
        RECT 2394.860 147.940 2395.120 148.200 ;
      LAYER met2 ;
        RECT 602.490 500.000 602.770 504.000 ;
        RECT 602.530 499.790 602.670 500.000 ;
        RECT 602.470 499.470 602.730 499.790 ;
        RECT 602.700 498.450 602.960 498.770 ;
        RECT 602.760 148.230 602.900 498.450 ;
        RECT 602.700 147.910 602.960 148.230 ;
        RECT 2394.860 147.910 2395.120 148.230 ;
        RECT 2394.920 82.870 2395.060 147.910 ;
        RECT 2394.920 82.730 2395.520 82.870 ;
        RECT 2395.380 2.400 2395.520 82.730 ;
        RECT 2395.170 -4.800 2395.730 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 603.130 168.880 603.450 168.940 ;
        RECT 2408.170 168.880 2408.490 168.940 ;
        RECT 603.130 168.740 2408.490 168.880 ;
        RECT 603.130 168.680 603.450 168.740 ;
        RECT 2408.170 168.680 2408.490 168.740 ;
      LAYER via ;
        RECT 603.160 168.680 603.420 168.940 ;
        RECT 2408.200 168.680 2408.460 168.940 ;
      LAYER met2 ;
        RECT 603.870 500.000 604.150 504.000 ;
        RECT 603.910 499.815 604.050 500.000 ;
        RECT 603.840 499.445 604.120 499.815 ;
        RECT 603.150 484.315 603.430 484.685 ;
        RECT 603.220 168.970 603.360 484.315 ;
        RECT 603.160 168.650 603.420 168.970 ;
        RECT 2408.200 168.650 2408.460 168.970 ;
        RECT 2408.260 82.870 2408.400 168.650 ;
        RECT 2408.260 82.730 2412.080 82.870 ;
        RECT 2411.940 2.400 2412.080 82.730 ;
        RECT 2411.730 -4.800 2412.290 2.400 ;
      LAYER via2 ;
        RECT 603.840 499.490 604.120 499.770 ;
        RECT 603.150 484.360 603.430 484.640 ;
      LAYER met3 ;
        RECT 603.815 499.620 604.145 499.795 ;
        RECT 603.790 499.610 604.170 499.620 ;
        RECT 603.790 499.310 604.430 499.610 ;
        RECT 603.790 499.300 604.170 499.310 ;
        RECT 603.790 485.330 604.170 485.340 ;
        RECT 602.910 485.030 604.170 485.330 ;
        RECT 602.910 484.665 603.210 485.030 ;
        RECT 603.790 485.020 604.170 485.030 ;
        RECT 602.910 484.350 603.455 484.665 ;
        RECT 603.125 484.335 603.455 484.350 ;
      LAYER via3 ;
        RECT 603.820 499.300 604.140 499.620 ;
        RECT 603.820 485.020 604.140 485.340 ;
      LAYER met4 ;
        RECT 603.815 499.295 604.145 499.625 ;
        RECT 603.830 485.345 604.130 499.295 ;
        RECT 603.815 485.015 604.145 485.345 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2421.970 17.920 2422.290 17.980 ;
        RECT 2428.410 17.920 2428.730 17.980 ;
        RECT 2421.970 17.780 2428.730 17.920 ;
        RECT 2421.970 17.720 2422.290 17.780 ;
        RECT 2428.410 17.720 2428.730 17.780 ;
      LAYER via ;
        RECT 2422.000 17.720 2422.260 17.980 ;
        RECT 2428.440 17.720 2428.700 17.980 ;
      LAYER met2 ;
        RECT 605.250 500.000 605.530 504.000 ;
        RECT 605.290 499.815 605.430 500.000 ;
        RECT 605.220 499.445 605.500 499.815 ;
        RECT 2421.990 175.595 2422.270 175.965 ;
        RECT 2422.060 18.010 2422.200 175.595 ;
        RECT 2422.000 17.690 2422.260 18.010 ;
        RECT 2428.440 17.690 2428.700 18.010 ;
        RECT 2428.500 2.400 2428.640 17.690 ;
        RECT 2428.290 -4.800 2428.850 2.400 ;
      LAYER via2 ;
        RECT 605.220 499.490 605.500 499.770 ;
        RECT 2421.990 175.640 2422.270 175.920 ;
      LAYER met3 ;
        RECT 605.195 499.780 605.525 499.795 ;
        RECT 604.980 499.465 605.525 499.780 ;
        RECT 604.980 498.940 605.280 499.465 ;
        RECT 604.710 498.630 605.280 498.940 ;
        RECT 604.710 498.620 605.090 498.630 ;
        RECT 604.710 175.930 605.090 175.940 ;
        RECT 2421.965 175.930 2422.295 175.945 ;
        RECT 604.710 175.630 2422.295 175.930 ;
        RECT 604.710 175.620 605.090 175.630 ;
        RECT 2421.965 175.615 2422.295 175.630 ;
      LAYER via3 ;
        RECT 604.740 498.620 605.060 498.940 ;
        RECT 604.740 175.620 605.060 175.940 ;
      LAYER met4 ;
        RECT 604.735 498.615 605.065 498.945 ;
        RECT 604.750 175.945 605.050 498.615 ;
        RECT 604.735 175.615 605.065 175.945 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.580 500.180 606.900 500.440 ;
        RECT 606.670 498.340 606.810 500.180 ;
        RECT 607.730 498.340 608.050 498.400 ;
        RECT 606.670 498.200 608.050 498.340 ;
        RECT 607.730 498.140 608.050 498.200 ;
      LAYER via ;
        RECT 606.610 500.180 606.870 500.440 ;
        RECT 607.760 498.140 608.020 498.400 ;
      LAYER met2 ;
        RECT 606.630 500.470 606.910 504.000 ;
        RECT 606.610 500.150 606.910 500.470 ;
        RECT 606.630 500.000 606.910 500.150 ;
        RECT 607.760 498.110 608.020 498.430 ;
        RECT 607.820 479.925 607.960 498.110 ;
        RECT 607.750 479.555 608.030 479.925 ;
        RECT 2442.690 479.555 2442.970 479.925 ;
        RECT 2442.760 82.870 2442.900 479.555 ;
        RECT 2442.760 82.730 2445.200 82.870 ;
        RECT 2445.060 2.400 2445.200 82.730 ;
        RECT 2444.850 -4.800 2445.410 2.400 ;
      LAYER via2 ;
        RECT 607.750 479.600 608.030 479.880 ;
        RECT 2442.690 479.600 2442.970 479.880 ;
      LAYER met3 ;
        RECT 607.725 479.890 608.055 479.905 ;
        RECT 2442.665 479.890 2442.995 479.905 ;
        RECT 607.725 479.590 2442.995 479.890 ;
        RECT 607.725 479.575 608.055 479.590 ;
        RECT 2442.665 479.575 2442.995 479.590 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.960 500.720 608.280 500.780 ;
        RECT 605.520 500.580 608.280 500.720 ;
        RECT 605.520 498.000 605.660 500.580 ;
        RECT 607.960 500.520 608.280 500.580 ;
        RECT 607.270 498.000 607.590 498.060 ;
        RECT 605.520 497.860 607.590 498.000 ;
        RECT 607.270 497.800 607.590 497.860 ;
        RECT 607.270 475.900 607.590 475.960 ;
        RECT 609.110 475.900 609.430 475.960 ;
        RECT 607.270 475.760 609.430 475.900 ;
        RECT 607.270 475.700 607.590 475.760 ;
        RECT 609.110 475.700 609.430 475.760 ;
        RECT 609.110 86.600 609.430 86.660 ;
        RECT 2456.470 86.600 2456.790 86.660 ;
        RECT 609.110 86.460 2456.790 86.600 ;
        RECT 609.110 86.400 609.430 86.460 ;
        RECT 2456.470 86.400 2456.790 86.460 ;
      LAYER via ;
        RECT 607.990 500.520 608.250 500.780 ;
        RECT 607.300 497.800 607.560 498.060 ;
        RECT 607.300 475.700 607.560 475.960 ;
        RECT 609.140 475.700 609.400 475.960 ;
        RECT 609.140 86.400 609.400 86.660 ;
        RECT 2456.500 86.400 2456.760 86.660 ;
      LAYER met2 ;
        RECT 608.010 500.810 608.290 504.000 ;
        RECT 607.990 500.490 608.290 500.810 ;
        RECT 608.010 500.000 608.290 500.490 ;
        RECT 607.300 497.770 607.560 498.090 ;
        RECT 607.360 475.990 607.500 497.770 ;
        RECT 607.300 475.670 607.560 475.990 ;
        RECT 609.140 475.670 609.400 475.990 ;
        RECT 609.200 86.690 609.340 475.670 ;
        RECT 609.140 86.370 609.400 86.690 ;
        RECT 2456.500 86.370 2456.760 86.690 ;
        RECT 2456.560 82.870 2456.700 86.370 ;
        RECT 2456.560 82.730 2461.760 82.870 ;
        RECT 2461.620 2.400 2461.760 82.730 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 609.340 499.360 609.660 499.420 ;
        RECT 608.740 499.220 609.660 499.360 ;
        RECT 608.740 497.720 608.880 499.220 ;
        RECT 609.340 499.160 609.660 499.220 ;
        RECT 608.650 497.460 608.970 497.720 ;
        RECT 608.650 86.260 608.970 86.320 ;
        RECT 2477.630 86.260 2477.950 86.320 ;
        RECT 608.650 86.120 2477.950 86.260 ;
        RECT 608.650 86.060 608.970 86.120 ;
        RECT 2477.630 86.060 2477.950 86.120 ;
      LAYER via ;
        RECT 609.370 499.160 609.630 499.420 ;
        RECT 608.680 497.460 608.940 497.720 ;
        RECT 608.680 86.060 608.940 86.320 ;
        RECT 2477.660 86.060 2477.920 86.320 ;
      LAYER met2 ;
        RECT 609.390 500.000 609.670 504.000 ;
        RECT 609.430 499.450 609.570 500.000 ;
        RECT 609.370 499.130 609.630 499.450 ;
        RECT 608.680 497.430 608.940 497.750 ;
        RECT 608.740 86.350 608.880 497.430 ;
        RECT 608.680 86.030 608.940 86.350 ;
        RECT 2477.660 86.030 2477.920 86.350 ;
        RECT 2477.720 82.870 2477.860 86.030 ;
        RECT 2477.720 82.730 2478.320 82.870 ;
        RECT 2478.180 2.400 2478.320 82.730 ;
        RECT 2477.970 -4.800 2478.530 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 610.030 480.660 610.350 480.720 ;
        RECT 2490.970 480.660 2491.290 480.720 ;
        RECT 610.030 480.520 2491.290 480.660 ;
        RECT 610.030 480.460 610.350 480.520 ;
        RECT 2490.970 480.460 2491.290 480.520 ;
      LAYER via ;
        RECT 610.060 480.460 610.320 480.720 ;
        RECT 2491.000 480.460 2491.260 480.720 ;
      LAYER met2 ;
        RECT 610.770 500.000 611.050 504.000 ;
        RECT 610.810 498.680 610.950 500.000 ;
        RECT 610.580 498.540 610.950 498.680 ;
        RECT 610.580 498.000 610.720 498.540 ;
        RECT 610.120 497.860 610.720 498.000 ;
        RECT 610.120 480.750 610.260 497.860 ;
        RECT 610.060 480.430 610.320 480.750 ;
        RECT 2491.000 480.430 2491.260 480.750 ;
        RECT 2491.060 82.870 2491.200 480.430 ;
        RECT 2491.060 82.730 2494.880 82.870 ;
        RECT 2494.740 2.400 2494.880 82.730 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2505.230 17.920 2505.550 17.980 ;
        RECT 2511.210 17.920 2511.530 17.980 ;
        RECT 2505.230 17.780 2511.530 17.920 ;
        RECT 2505.230 17.720 2505.550 17.780 ;
        RECT 2511.210 17.720 2511.530 17.780 ;
      LAYER via ;
        RECT 2505.260 17.720 2505.520 17.980 ;
        RECT 2511.240 17.720 2511.500 17.980 ;
      LAYER met2 ;
        RECT 612.150 500.000 612.430 504.000 ;
        RECT 612.190 498.965 612.330 500.000 ;
        RECT 612.120 498.595 612.400 498.965 ;
        RECT 2505.250 85.835 2505.530 86.205 ;
        RECT 2505.320 18.010 2505.460 85.835 ;
        RECT 2505.260 17.690 2505.520 18.010 ;
        RECT 2511.240 17.690 2511.500 18.010 ;
        RECT 2511.300 2.400 2511.440 17.690 ;
        RECT 2511.090 -4.800 2511.650 2.400 ;
      LAYER via2 ;
        RECT 612.120 498.640 612.400 498.920 ;
        RECT 2505.250 85.880 2505.530 86.160 ;
      LAYER met3 ;
        RECT 612.095 498.940 612.425 498.945 ;
        RECT 612.070 498.930 612.450 498.940 ;
        RECT 611.640 498.630 612.450 498.930 ;
        RECT 612.070 498.620 612.450 498.630 ;
        RECT 612.095 498.615 612.425 498.620 ;
        RECT 612.070 86.170 612.450 86.180 ;
        RECT 2505.225 86.170 2505.555 86.185 ;
        RECT 612.070 85.870 2505.555 86.170 ;
        RECT 612.070 85.860 612.450 85.870 ;
        RECT 2505.225 85.855 2505.555 85.870 ;
      LAYER via3 ;
        RECT 612.100 498.620 612.420 498.940 ;
        RECT 612.100 85.860 612.420 86.180 ;
      LAYER met4 ;
        RECT 612.095 498.615 612.425 498.945 ;
        RECT 612.110 86.185 612.410 498.615 ;
        RECT 612.095 85.855 612.425 86.185 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 475.480 499.360 475.800 499.420 ;
        RECT 475.480 499.220 478.240 499.360 ;
        RECT 475.480 499.160 475.800 499.220 ;
        RECT 475.710 497.320 476.030 497.380 ;
        RECT 478.100 497.320 478.240 499.220 ;
        RECT 475.710 497.180 478.240 497.320 ;
        RECT 475.710 497.120 476.030 497.180 ;
      LAYER via ;
        RECT 475.510 499.160 475.770 499.420 ;
        RECT 475.740 497.120 476.000 497.380 ;
      LAYER met2 ;
        RECT 475.530 500.000 475.810 504.000 ;
        RECT 475.570 499.450 475.710 500.000 ;
        RECT 475.510 499.130 475.770 499.450 ;
        RECT 475.740 497.090 476.000 497.410 ;
        RECT 475.800 489.445 475.940 497.090 ;
        RECT 475.730 489.075 476.010 489.445 ;
        RECT 869.490 181.715 869.770 182.085 ;
        RECT 869.560 82.870 869.700 181.715 ;
        RECT 869.560 82.730 872.000 82.870 ;
        RECT 871.860 2.400 872.000 82.730 ;
        RECT 871.650 -4.800 872.210 2.400 ;
      LAYER via2 ;
        RECT 475.730 489.120 476.010 489.400 ;
        RECT 869.490 181.760 869.770 182.040 ;
      LAYER met3 ;
        RECT 474.070 489.410 474.450 489.420 ;
        RECT 475.705 489.410 476.035 489.425 ;
        RECT 474.070 489.110 476.035 489.410 ;
        RECT 474.070 489.100 474.450 489.110 ;
        RECT 475.705 489.095 476.035 489.110 ;
        RECT 474.070 182.050 474.450 182.060 ;
        RECT 869.465 182.050 869.795 182.065 ;
        RECT 474.070 181.750 869.795 182.050 ;
        RECT 474.070 181.740 474.450 181.750 ;
        RECT 869.465 181.735 869.795 181.750 ;
      LAYER via3 ;
        RECT 474.100 489.100 474.420 489.420 ;
        RECT 474.100 181.740 474.420 182.060 ;
      LAYER met4 ;
        RECT 474.095 489.095 474.425 489.425 ;
        RECT 474.110 182.065 474.410 489.095 ;
        RECT 474.095 181.735 474.425 182.065 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.480 499.500 613.800 499.760 ;
        RECT 613.570 497.720 613.710 499.500 ;
        RECT 613.250 497.520 613.710 497.720 ;
        RECT 613.250 497.460 613.570 497.520 ;
      LAYER via ;
        RECT 613.510 499.500 613.770 499.760 ;
        RECT 613.280 497.460 613.540 497.720 ;
      LAYER met2 ;
        RECT 613.530 500.000 613.810 504.000 ;
        RECT 613.570 499.790 613.710 500.000 ;
        RECT 613.510 499.470 613.770 499.790 ;
        RECT 613.280 497.430 613.540 497.750 ;
        RECT 613.340 484.005 613.480 497.430 ;
        RECT 613.270 483.635 613.550 484.005 ;
        RECT 2525.490 93.315 2525.770 93.685 ;
        RECT 2525.560 82.870 2525.700 93.315 ;
        RECT 2525.560 82.730 2528.000 82.870 ;
        RECT 2527.860 2.400 2528.000 82.730 ;
        RECT 2527.650 -4.800 2528.210 2.400 ;
      LAYER via2 ;
        RECT 613.270 483.680 613.550 483.960 ;
        RECT 2525.490 93.360 2525.770 93.640 ;
      LAYER met3 ;
        RECT 611.150 483.970 611.530 483.980 ;
        RECT 613.245 483.970 613.575 483.985 ;
        RECT 611.150 483.670 613.575 483.970 ;
        RECT 611.150 483.660 611.530 483.670 ;
        RECT 613.245 483.655 613.575 483.670 ;
        RECT 611.150 93.650 611.530 93.660 ;
        RECT 2525.465 93.650 2525.795 93.665 ;
        RECT 611.150 93.350 2525.795 93.650 ;
        RECT 611.150 93.340 611.530 93.350 ;
        RECT 2525.465 93.335 2525.795 93.350 ;
      LAYER via3 ;
        RECT 611.180 483.660 611.500 483.980 ;
        RECT 611.180 93.340 611.500 93.660 ;
      LAYER met4 ;
        RECT 611.175 483.655 611.505 483.985 ;
        RECT 611.190 93.665 611.490 483.655 ;
        RECT 611.175 93.335 611.505 93.665 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 471.820 615.410 471.880 ;
        RECT 616.930 471.820 617.250 471.880 ;
        RECT 615.090 471.680 617.250 471.820 ;
        RECT 615.090 471.620 615.410 471.680 ;
        RECT 616.930 471.620 617.250 471.680 ;
        RECT 616.930 403.480 617.250 403.540 ;
        RECT 2539.270 403.480 2539.590 403.540 ;
        RECT 616.930 403.340 2539.590 403.480 ;
        RECT 616.930 403.280 617.250 403.340 ;
        RECT 2539.270 403.280 2539.590 403.340 ;
      LAYER via ;
        RECT 615.120 471.620 615.380 471.880 ;
        RECT 616.960 471.620 617.220 471.880 ;
        RECT 616.960 403.280 617.220 403.540 ;
        RECT 2539.300 403.280 2539.560 403.540 ;
      LAYER met2 ;
        RECT 614.910 500.000 615.190 504.000 ;
        RECT 614.950 498.850 615.090 500.000 ;
        RECT 614.950 498.710 615.320 498.850 ;
        RECT 615.180 471.910 615.320 498.710 ;
        RECT 615.120 471.590 615.380 471.910 ;
        RECT 616.960 471.590 617.220 471.910 ;
        RECT 617.020 403.570 617.160 471.590 ;
        RECT 616.960 403.250 617.220 403.570 ;
        RECT 2539.300 403.250 2539.560 403.570 ;
        RECT 2539.360 82.870 2539.500 403.250 ;
        RECT 2539.360 82.730 2544.560 82.870 ;
        RECT 2544.420 2.400 2544.560 82.730 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 616.240 499.500 616.560 499.760 ;
        RECT 616.330 498.400 616.470 499.500 ;
        RECT 616.330 498.200 616.790 498.400 ;
        RECT 616.470 498.140 616.790 498.200 ;
        RECT 616.470 474.880 616.790 474.940 ;
        RECT 617.390 474.880 617.710 474.940 ;
        RECT 616.470 474.740 617.710 474.880 ;
        RECT 616.470 474.680 616.790 474.740 ;
        RECT 617.390 474.680 617.710 474.740 ;
        RECT 617.390 410.620 617.710 410.680 ;
        RECT 2560.430 410.620 2560.750 410.680 ;
        RECT 617.390 410.480 2560.750 410.620 ;
        RECT 617.390 410.420 617.710 410.480 ;
        RECT 2560.430 410.420 2560.750 410.480 ;
      LAYER via ;
        RECT 616.270 499.500 616.530 499.760 ;
        RECT 616.500 498.140 616.760 498.400 ;
        RECT 616.500 474.680 616.760 474.940 ;
        RECT 617.420 474.680 617.680 474.940 ;
        RECT 617.420 410.420 617.680 410.680 ;
        RECT 2560.460 410.420 2560.720 410.680 ;
      LAYER met2 ;
        RECT 616.290 500.000 616.570 504.000 ;
        RECT 616.330 499.790 616.470 500.000 ;
        RECT 616.270 499.470 616.530 499.790 ;
        RECT 616.500 498.110 616.760 498.430 ;
        RECT 616.560 474.970 616.700 498.110 ;
        RECT 616.500 474.650 616.760 474.970 ;
        RECT 617.420 474.650 617.680 474.970 ;
        RECT 617.480 410.710 617.620 474.650 ;
        RECT 617.420 410.390 617.680 410.710 ;
        RECT 2560.460 410.390 2560.720 410.710 ;
        RECT 2560.520 82.870 2560.660 410.390 ;
        RECT 2560.520 82.730 2561.120 82.870 ;
        RECT 2560.980 2.400 2561.120 82.730 ;
        RECT 2560.770 -4.800 2561.330 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.620 499.700 617.940 499.760 ;
        RECT 617.620 499.560 619.230 499.700 ;
        RECT 617.620 499.500 617.940 499.560 ;
        RECT 619.090 498.400 619.230 499.560 ;
        RECT 619.090 498.200 619.550 498.400 ;
        RECT 619.230 498.140 619.550 498.200 ;
        RECT 619.230 480.320 619.550 480.380 ;
        RECT 2573.770 480.320 2574.090 480.380 ;
        RECT 619.230 480.180 2574.090 480.320 ;
        RECT 619.230 480.120 619.550 480.180 ;
        RECT 2573.770 480.120 2574.090 480.180 ;
      LAYER via ;
        RECT 617.650 499.500 617.910 499.760 ;
        RECT 619.260 498.140 619.520 498.400 ;
        RECT 619.260 480.120 619.520 480.380 ;
        RECT 2573.800 480.120 2574.060 480.380 ;
      LAYER met2 ;
        RECT 617.670 500.000 617.950 504.000 ;
        RECT 617.710 499.790 617.850 500.000 ;
        RECT 617.650 499.470 617.910 499.790 ;
        RECT 619.260 498.110 619.520 498.430 ;
        RECT 619.320 480.410 619.460 498.110 ;
        RECT 619.260 480.090 619.520 480.410 ;
        RECT 2573.800 480.090 2574.060 480.410 ;
        RECT 2573.860 82.870 2574.000 480.090 ;
        RECT 2573.860 82.730 2577.680 82.870 ;
        RECT 2577.540 2.400 2577.680 82.730 ;
        RECT 2577.330 -4.800 2577.890 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 471.140 615.410 471.200 ;
        RECT 618.770 471.140 619.090 471.200 ;
        RECT 615.090 471.000 619.090 471.140 ;
        RECT 615.090 470.940 615.410 471.000 ;
        RECT 618.770 470.940 619.090 471.000 ;
        RECT 615.090 93.400 615.410 93.460 ;
        RECT 2587.570 93.400 2587.890 93.460 ;
        RECT 615.090 93.260 2587.890 93.400 ;
        RECT 615.090 93.200 615.410 93.260 ;
        RECT 2587.570 93.200 2587.890 93.260 ;
        RECT 2587.570 37.640 2587.890 37.700 ;
        RECT 2594.010 37.640 2594.330 37.700 ;
        RECT 2587.570 37.500 2594.330 37.640 ;
        RECT 2587.570 37.440 2587.890 37.500 ;
        RECT 2594.010 37.440 2594.330 37.500 ;
      LAYER via ;
        RECT 615.120 470.940 615.380 471.200 ;
        RECT 618.800 470.940 619.060 471.200 ;
        RECT 615.120 93.200 615.380 93.460 ;
        RECT 2587.600 93.200 2587.860 93.460 ;
        RECT 2587.600 37.440 2587.860 37.700 ;
        RECT 2594.040 37.440 2594.300 37.700 ;
      LAYER met2 ;
        RECT 619.050 500.000 619.330 504.000 ;
        RECT 619.090 498.850 619.230 500.000 ;
        RECT 618.860 498.710 619.230 498.850 ;
        RECT 618.860 471.230 619.000 498.710 ;
        RECT 615.120 470.910 615.380 471.230 ;
        RECT 618.800 470.910 619.060 471.230 ;
        RECT 615.180 93.490 615.320 470.910 ;
        RECT 615.120 93.170 615.380 93.490 ;
        RECT 2587.600 93.170 2587.860 93.490 ;
        RECT 2587.660 37.730 2587.800 93.170 ;
        RECT 2587.600 37.410 2587.860 37.730 ;
        RECT 2594.040 37.410 2594.300 37.730 ;
        RECT 2594.100 2.400 2594.240 37.410 ;
        RECT 2593.890 -4.800 2594.450 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 620.380 499.500 620.700 499.760 ;
        RECT 620.470 498.740 620.610 499.500 ;
        RECT 620.150 498.540 620.610 498.740 ;
        RECT 620.150 498.480 620.470 498.540 ;
      LAYER via ;
        RECT 620.410 499.500 620.670 499.760 ;
        RECT 620.180 498.480 620.440 498.740 ;
      LAYER met2 ;
        RECT 620.430 500.000 620.710 504.000 ;
        RECT 620.470 499.790 620.610 500.000 ;
        RECT 620.410 499.470 620.670 499.790 ;
        RECT 620.180 498.450 620.440 498.770 ;
        RECT 620.240 491.485 620.380 498.450 ;
        RECT 620.170 491.115 620.450 491.485 ;
        RECT 2608.290 478.875 2608.570 479.245 ;
        RECT 2608.360 82.870 2608.500 478.875 ;
        RECT 2608.360 82.730 2610.800 82.870 ;
        RECT 2610.660 2.400 2610.800 82.730 ;
        RECT 2610.450 -4.800 2611.010 2.400 ;
      LAYER via2 ;
        RECT 620.170 491.160 620.450 491.440 ;
        RECT 2608.290 478.920 2608.570 479.200 ;
      LAYER met3 ;
        RECT 613.910 491.450 614.290 491.460 ;
        RECT 620.145 491.450 620.475 491.465 ;
        RECT 613.910 491.150 620.475 491.450 ;
        RECT 613.910 491.140 614.290 491.150 ;
        RECT 620.145 491.135 620.475 491.150 ;
        RECT 613.910 479.210 614.290 479.220 ;
        RECT 2608.265 479.210 2608.595 479.225 ;
        RECT 613.910 478.910 2608.595 479.210 ;
        RECT 613.910 478.900 614.290 478.910 ;
        RECT 2608.265 478.895 2608.595 478.910 ;
      LAYER via3 ;
        RECT 613.940 491.140 614.260 491.460 ;
        RECT 613.940 478.900 614.260 479.220 ;
      LAYER met4 ;
        RECT 613.935 491.135 614.265 491.465 ;
        RECT 613.950 479.225 614.250 491.135 ;
        RECT 613.935 478.895 614.265 479.225 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.760 499.360 622.080 499.420 ;
        RECT 621.760 499.220 623.600 499.360 ;
        RECT 621.760 499.160 622.080 499.220 ;
        RECT 623.460 499.080 623.600 499.220 ;
        RECT 623.370 498.820 623.690 499.080 ;
        RECT 623.370 93.060 623.690 93.120 ;
        RECT 2622.070 93.060 2622.390 93.120 ;
        RECT 623.370 92.920 2622.390 93.060 ;
        RECT 623.370 92.860 623.690 92.920 ;
        RECT 2622.070 92.860 2622.390 92.920 ;
      LAYER via ;
        RECT 621.790 499.160 622.050 499.420 ;
        RECT 623.400 498.820 623.660 499.080 ;
        RECT 623.400 92.860 623.660 93.120 ;
        RECT 2622.100 92.860 2622.360 93.120 ;
      LAYER met2 ;
        RECT 621.810 500.000 622.090 504.000 ;
        RECT 621.850 499.450 621.990 500.000 ;
        RECT 621.790 499.130 622.050 499.450 ;
        RECT 623.400 498.790 623.660 499.110 ;
        RECT 623.460 93.150 623.600 498.790 ;
        RECT 623.400 92.830 623.660 93.150 ;
        RECT 2622.100 92.830 2622.360 93.150 ;
        RECT 2622.160 82.870 2622.300 92.830 ;
        RECT 2622.160 82.730 2627.360 82.870 ;
        RECT 2627.220 2.400 2627.360 82.730 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.510 479.980 627.830 480.040 ;
        RECT 2642.770 479.980 2643.090 480.040 ;
        RECT 627.510 479.840 2643.090 479.980 ;
        RECT 627.510 479.780 627.830 479.840 ;
        RECT 2642.770 479.780 2643.090 479.840 ;
      LAYER via ;
        RECT 627.540 479.780 627.800 480.040 ;
        RECT 2642.800 479.780 2643.060 480.040 ;
      LAYER met2 ;
        RECT 623.190 500.000 623.470 504.000 ;
        RECT 623.230 499.645 623.370 500.000 ;
        RECT 623.160 499.275 623.440 499.645 ;
        RECT 627.530 497.235 627.810 497.605 ;
        RECT 627.600 480.070 627.740 497.235 ;
        RECT 627.540 479.750 627.800 480.070 ;
        RECT 2642.800 479.750 2643.060 480.070 ;
        RECT 2642.860 82.870 2643.000 479.750 ;
        RECT 2642.860 82.730 2643.920 82.870 ;
        RECT 2643.780 2.400 2643.920 82.730 ;
        RECT 2643.570 -4.800 2644.130 2.400 ;
      LAYER via2 ;
        RECT 623.160 499.320 623.440 499.600 ;
        RECT 627.530 497.280 627.810 497.560 ;
      LAYER met3 ;
        RECT 623.135 499.295 623.465 499.625 ;
        RECT 623.150 497.570 623.450 499.295 ;
        RECT 627.505 497.570 627.835 497.585 ;
        RECT 623.150 497.270 627.835 497.570 ;
        RECT 627.505 497.255 627.835 497.270 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 624.290 176.020 624.610 176.080 ;
        RECT 2656.570 176.020 2656.890 176.080 ;
        RECT 624.290 175.880 2656.890 176.020 ;
        RECT 624.290 175.820 624.610 175.880 ;
        RECT 2656.570 175.820 2656.890 175.880 ;
      LAYER via ;
        RECT 624.320 175.820 624.580 176.080 ;
        RECT 2656.600 175.820 2656.860 176.080 ;
      LAYER met2 ;
        RECT 624.570 500.000 624.850 504.000 ;
        RECT 624.610 499.020 624.750 500.000 ;
        RECT 624.380 498.880 624.750 499.020 ;
        RECT 624.380 176.110 624.520 498.880 ;
        RECT 624.320 175.790 624.580 176.110 ;
        RECT 2656.600 175.790 2656.860 176.110 ;
        RECT 2656.660 82.870 2656.800 175.790 ;
        RECT 2656.660 82.730 2660.480 82.870 ;
        RECT 2660.340 2.400 2660.480 82.730 ;
        RECT 2660.130 -4.800 2660.690 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2670.370 3.640 2670.690 3.700 ;
        RECT 2676.810 3.640 2677.130 3.700 ;
        RECT 2670.370 3.500 2677.130 3.640 ;
        RECT 2670.370 3.440 2670.690 3.500 ;
        RECT 2676.810 3.440 2677.130 3.500 ;
      LAYER via ;
        RECT 2670.400 3.440 2670.660 3.700 ;
        RECT 2676.840 3.440 2677.100 3.700 ;
      LAYER met2 ;
        RECT 625.950 500.000 626.230 504.000 ;
        RECT 625.990 498.850 626.130 500.000 ;
        RECT 625.990 498.710 626.360 498.850 ;
        RECT 626.220 484.005 626.360 498.710 ;
        RECT 626.150 483.635 626.430 484.005 ;
        RECT 2670.390 92.635 2670.670 93.005 ;
        RECT 2670.460 3.730 2670.600 92.635 ;
        RECT 2670.400 3.410 2670.660 3.730 ;
        RECT 2676.840 3.410 2677.100 3.730 ;
        RECT 2676.900 2.400 2677.040 3.410 ;
        RECT 2676.690 -4.800 2677.250 2.400 ;
      LAYER via2 ;
        RECT 626.150 483.680 626.430 483.960 ;
        RECT 2670.390 92.680 2670.670 92.960 ;
      LAYER met3 ;
        RECT 626.125 483.970 626.455 483.985 ;
        RECT 626.790 483.970 627.170 483.980 ;
        RECT 626.125 483.670 627.170 483.970 ;
        RECT 626.125 483.655 626.455 483.670 ;
        RECT 626.790 483.660 627.170 483.670 ;
        RECT 626.790 92.970 627.170 92.980 ;
        RECT 2670.365 92.970 2670.695 92.985 ;
        RECT 626.790 92.670 2670.695 92.970 ;
        RECT 626.790 92.660 627.170 92.670 ;
        RECT 2670.365 92.655 2670.695 92.670 ;
      LAYER via3 ;
        RECT 626.820 483.660 627.140 483.980 ;
        RECT 626.820 92.660 627.140 92.980 ;
      LAYER met4 ;
        RECT 626.815 483.655 627.145 483.985 ;
        RECT 626.830 92.985 627.130 483.655 ;
        RECT 626.815 92.655 627.145 92.985 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 481.680 476.490 481.740 ;
        RECT 883.270 481.680 883.590 481.740 ;
        RECT 476.170 481.540 883.590 481.680 ;
        RECT 476.170 481.480 476.490 481.540 ;
        RECT 883.270 481.480 883.590 481.540 ;
      LAYER via ;
        RECT 476.200 481.480 476.460 481.740 ;
        RECT 883.300 481.480 883.560 481.740 ;
      LAYER met2 ;
        RECT 476.910 500.000 477.190 504.000 ;
        RECT 476.950 499.020 477.090 500.000 ;
        RECT 476.950 498.880 477.320 499.020 ;
        RECT 477.180 497.320 477.320 498.880 ;
        RECT 476.720 497.180 477.320 497.320 ;
        RECT 476.720 491.880 476.860 497.180 ;
        RECT 476.260 491.740 476.860 491.880 ;
        RECT 476.260 481.770 476.400 491.740 ;
        RECT 476.200 481.450 476.460 481.770 ;
        RECT 883.300 481.450 883.560 481.770 ;
        RECT 883.360 82.870 883.500 481.450 ;
        RECT 883.360 82.730 888.560 82.870 ;
        RECT 888.420 2.400 888.560 82.730 ;
        RECT 888.210 -4.800 888.770 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.330 500.000 627.610 504.000 ;
        RECT 627.370 498.340 627.510 500.000 ;
        RECT 627.140 498.200 627.510 498.340 ;
        RECT 627.140 485.365 627.280 498.200 ;
        RECT 627.070 484.995 627.350 485.365 ;
        RECT 2691.090 183.075 2691.370 183.445 ;
        RECT 2691.160 82.870 2691.300 183.075 ;
        RECT 2691.160 82.730 2693.600 82.870 ;
        RECT 2693.460 2.400 2693.600 82.730 ;
        RECT 2693.250 -4.800 2693.810 2.400 ;
      LAYER via2 ;
        RECT 627.070 485.040 627.350 485.320 ;
        RECT 2691.090 183.120 2691.370 183.400 ;
      LAYER met3 ;
        RECT 624.950 485.330 625.330 485.340 ;
        RECT 627.045 485.330 627.375 485.345 ;
        RECT 624.950 485.030 627.375 485.330 ;
        RECT 624.950 485.020 625.330 485.030 ;
        RECT 627.045 485.015 627.375 485.030 ;
        RECT 624.950 183.410 625.330 183.420 ;
        RECT 2691.065 183.410 2691.395 183.425 ;
        RECT 624.950 183.110 2691.395 183.410 ;
        RECT 624.950 183.100 625.330 183.110 ;
        RECT 2691.065 183.095 2691.395 183.110 ;
      LAYER via3 ;
        RECT 624.980 485.020 625.300 485.340 ;
        RECT 624.980 183.100 625.300 183.420 ;
      LAYER met4 ;
        RECT 624.975 485.015 625.305 485.345 ;
        RECT 624.990 183.425 625.290 485.015 ;
        RECT 624.975 183.095 625.305 183.425 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.660 500.180 628.980 500.440 ;
        RECT 628.750 500.040 628.890 500.180 ;
        RECT 628.750 499.900 629.810 500.040 ;
        RECT 629.670 498.060 629.810 499.900 ;
        RECT 629.670 497.860 630.130 498.060 ;
        RECT 629.810 497.800 630.130 497.860 ;
        RECT 629.810 79.800 630.130 79.860 ;
        RECT 2709.930 79.800 2710.250 79.860 ;
        RECT 629.810 79.660 2710.250 79.800 ;
        RECT 629.810 79.600 630.130 79.660 ;
        RECT 2709.930 79.600 2710.250 79.660 ;
      LAYER via ;
        RECT 628.690 500.180 628.950 500.440 ;
        RECT 629.840 497.800 630.100 498.060 ;
        RECT 629.840 79.600 630.100 79.860 ;
        RECT 2709.960 79.600 2710.220 79.860 ;
      LAYER met2 ;
        RECT 628.710 500.470 628.990 504.000 ;
        RECT 628.690 500.150 628.990 500.470 ;
        RECT 628.710 500.000 628.990 500.150 ;
        RECT 629.840 497.770 630.100 498.090 ;
        RECT 629.900 79.890 630.040 497.770 ;
        RECT 629.840 79.570 630.100 79.890 ;
        RECT 2709.960 79.570 2710.220 79.890 ;
        RECT 2710.020 2.400 2710.160 79.570 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 630.040 499.500 630.360 499.760 ;
        RECT 630.130 498.340 630.270 499.500 ;
        RECT 630.130 498.200 631.880 498.340 ;
        RECT 631.740 497.660 631.880 498.200 ;
        RECT 632.570 497.660 632.890 497.720 ;
        RECT 631.740 497.520 632.890 497.660 ;
        RECT 632.570 497.460 632.890 497.520 ;
        RECT 632.570 479.640 632.890 479.700 ;
        RECT 2725.570 479.640 2725.890 479.700 ;
        RECT 632.570 479.500 2725.890 479.640 ;
        RECT 632.570 479.440 632.890 479.500 ;
        RECT 2725.570 479.440 2725.890 479.500 ;
      LAYER via ;
        RECT 630.070 499.500 630.330 499.760 ;
        RECT 632.600 497.460 632.860 497.720 ;
        RECT 632.600 479.440 632.860 479.700 ;
        RECT 2725.600 479.440 2725.860 479.700 ;
      LAYER met2 ;
        RECT 630.090 500.000 630.370 504.000 ;
        RECT 630.130 499.790 630.270 500.000 ;
        RECT 630.070 499.470 630.330 499.790 ;
        RECT 632.600 497.430 632.860 497.750 ;
        RECT 632.660 479.730 632.800 497.430 ;
        RECT 632.600 479.410 632.860 479.730 ;
        RECT 2725.600 479.410 2725.860 479.730 ;
        RECT 2725.660 17.410 2725.800 479.410 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 631.420 499.500 631.740 499.760 ;
        RECT 631.510 498.740 631.650 499.500 ;
        RECT 631.190 498.540 631.650 498.740 ;
        RECT 631.190 498.480 631.510 498.540 ;
        RECT 2584.440 24.240 2608.270 24.380 ;
        RECT 627.970 24.040 628.290 24.100 ;
        RECT 2584.440 24.040 2584.580 24.240 ;
        RECT 627.970 23.900 2584.580 24.040 ;
        RECT 2608.130 24.040 2608.270 24.240 ;
        RECT 2743.050 24.040 2743.370 24.100 ;
        RECT 2608.130 23.900 2743.370 24.040 ;
        RECT 627.970 23.840 628.290 23.900 ;
        RECT 2743.050 23.840 2743.370 23.900 ;
      LAYER via ;
        RECT 631.450 499.500 631.710 499.760 ;
        RECT 631.220 498.480 631.480 498.740 ;
        RECT 628.000 23.840 628.260 24.100 ;
        RECT 2743.080 23.840 2743.340 24.100 ;
      LAYER met2 ;
        RECT 631.470 500.000 631.750 504.000 ;
        RECT 631.510 499.790 631.650 500.000 ;
        RECT 631.450 499.470 631.710 499.790 ;
        RECT 631.220 498.450 631.480 498.770 ;
        RECT 631.280 498.285 631.420 498.450 ;
        RECT 631.210 497.915 631.490 498.285 ;
        RECT 627.990 496.555 628.270 496.925 ;
        RECT 628.060 24.130 628.200 496.555 ;
        RECT 628.000 23.810 628.260 24.130 ;
        RECT 2743.080 23.810 2743.340 24.130 ;
        RECT 2743.140 2.400 2743.280 23.810 ;
        RECT 2742.930 -4.800 2743.490 2.400 ;
      LAYER via2 ;
        RECT 631.210 497.960 631.490 498.240 ;
        RECT 627.990 496.600 628.270 496.880 ;
      LAYER met3 ;
        RECT 631.185 498.250 631.515 498.265 ;
        RECT 630.510 497.950 631.515 498.250 ;
        RECT 627.965 496.890 628.295 496.905 ;
        RECT 630.510 496.890 630.810 497.950 ;
        RECT 631.185 497.935 631.515 497.950 ;
        RECT 627.965 496.590 630.810 496.890 ;
        RECT 627.965 496.575 628.295 496.590 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2753.630 17.920 2753.950 17.980 ;
        RECT 2759.610 17.920 2759.930 17.980 ;
        RECT 2753.630 17.780 2759.930 17.920 ;
        RECT 2753.630 17.720 2753.950 17.780 ;
        RECT 2759.610 17.720 2759.930 17.780 ;
      LAYER via ;
        RECT 2753.660 17.720 2753.920 17.980 ;
        RECT 2759.640 17.720 2759.900 17.980 ;
      LAYER met2 ;
        RECT 632.850 500.000 633.130 504.000 ;
        RECT 632.890 498.340 633.030 500.000 ;
        RECT 632.890 498.200 633.260 498.340 ;
        RECT 633.120 486.725 633.260 498.200 ;
        RECT 633.050 486.355 633.330 486.725 ;
        RECT 2753.650 99.435 2753.930 99.805 ;
        RECT 2753.720 18.010 2753.860 99.435 ;
        RECT 2753.660 17.690 2753.920 18.010 ;
        RECT 2759.640 17.690 2759.900 18.010 ;
        RECT 2759.700 2.400 2759.840 17.690 ;
        RECT 2759.490 -4.800 2760.050 2.400 ;
      LAYER via2 ;
        RECT 633.050 486.400 633.330 486.680 ;
        RECT 2753.650 99.480 2753.930 99.760 ;
      LAYER met3 ;
        RECT 633.025 486.690 633.355 486.705 ;
        RECT 634.150 486.690 634.530 486.700 ;
        RECT 633.025 486.390 634.530 486.690 ;
        RECT 633.025 486.375 633.355 486.390 ;
        RECT 634.150 486.380 634.530 486.390 ;
        RECT 634.150 99.770 634.530 99.780 ;
        RECT 2753.625 99.770 2753.955 99.785 ;
        RECT 634.150 99.470 2753.955 99.770 ;
        RECT 634.150 99.460 634.530 99.470 ;
        RECT 2753.625 99.455 2753.955 99.470 ;
      LAYER via3 ;
        RECT 634.180 486.380 634.500 486.700 ;
        RECT 634.180 99.460 634.500 99.780 ;
      LAYER met4 ;
        RECT 634.175 486.375 634.505 486.705 ;
        RECT 634.190 99.785 634.490 486.375 ;
        RECT 634.175 99.455 634.505 99.785 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.180 499.160 634.500 499.420 ;
        RECT 634.270 498.060 634.410 499.160 ;
        RECT 634.270 497.860 634.730 498.060 ;
        RECT 634.410 497.800 634.730 497.860 ;
      LAYER via ;
        RECT 634.210 499.160 634.470 499.420 ;
        RECT 634.440 497.800 634.700 498.060 ;
      LAYER met2 ;
        RECT 634.230 500.000 634.510 504.000 ;
        RECT 634.270 499.450 634.410 500.000 ;
        RECT 634.210 499.130 634.470 499.450 ;
        RECT 634.440 497.770 634.700 498.090 ;
        RECT 634.500 491.485 634.640 497.770 ;
        RECT 634.430 491.115 634.710 491.485 ;
        RECT 2773.890 182.395 2774.170 182.765 ;
        RECT 2773.960 82.870 2774.100 182.395 ;
        RECT 2773.960 82.730 2776.400 82.870 ;
        RECT 2776.260 2.400 2776.400 82.730 ;
        RECT 2776.050 -4.800 2776.610 2.400 ;
      LAYER via2 ;
        RECT 634.430 491.160 634.710 491.440 ;
        RECT 2773.890 182.440 2774.170 182.720 ;
      LAYER met3 ;
        RECT 632.310 491.450 632.690 491.460 ;
        RECT 634.405 491.450 634.735 491.465 ;
        RECT 632.310 491.150 634.735 491.450 ;
        RECT 632.310 491.140 632.690 491.150 ;
        RECT 634.405 491.135 634.735 491.150 ;
        RECT 632.310 182.730 632.690 182.740 ;
        RECT 2773.865 182.730 2774.195 182.745 ;
        RECT 632.310 182.430 2774.195 182.730 ;
        RECT 632.310 182.420 632.690 182.430 ;
        RECT 2773.865 182.415 2774.195 182.430 ;
      LAYER via3 ;
        RECT 632.340 491.140 632.660 491.460 ;
        RECT 632.340 182.420 632.660 182.740 ;
      LAYER met4 ;
        RECT 632.335 491.135 632.665 491.465 ;
        RECT 632.350 182.745 632.650 491.135 ;
        RECT 632.335 182.415 632.665 182.745 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.560 500.380 635.880 500.440 ;
        RECT 639.010 500.380 639.330 500.440 ;
        RECT 635.560 500.240 639.330 500.380 ;
        RECT 635.560 500.180 635.880 500.240 ;
        RECT 639.010 500.180 639.330 500.240 ;
        RECT 639.010 100.200 639.330 100.260 ;
        RECT 2787.670 100.200 2787.990 100.260 ;
        RECT 639.010 100.060 2787.990 100.200 ;
        RECT 639.010 100.000 639.330 100.060 ;
        RECT 2787.670 100.000 2787.990 100.060 ;
      LAYER via ;
        RECT 635.590 500.180 635.850 500.440 ;
        RECT 639.040 500.180 639.300 500.440 ;
        RECT 639.040 100.000 639.300 100.260 ;
        RECT 2787.700 100.000 2787.960 100.260 ;
      LAYER met2 ;
        RECT 635.610 500.470 635.890 504.000 ;
        RECT 635.590 500.150 635.890 500.470 ;
        RECT 639.040 500.150 639.300 500.470 ;
        RECT 635.610 500.000 635.890 500.150 ;
        RECT 639.100 100.290 639.240 500.150 ;
        RECT 639.040 99.970 639.300 100.290 ;
        RECT 2787.700 99.970 2787.960 100.290 ;
        RECT 2787.760 82.870 2787.900 99.970 ;
        RECT 2787.760 82.730 2792.960 82.870 ;
        RECT 2792.820 2.400 2792.960 82.730 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 637.170 99.860 637.490 99.920 ;
        RECT 2808.370 99.860 2808.690 99.920 ;
        RECT 637.170 99.720 2808.690 99.860 ;
        RECT 637.170 99.660 637.490 99.720 ;
        RECT 2808.370 99.660 2808.690 99.720 ;
      LAYER via ;
        RECT 637.200 99.660 637.460 99.920 ;
        RECT 2808.400 99.660 2808.660 99.920 ;
      LAYER met2 ;
        RECT 636.990 500.210 637.270 504.000 ;
        RECT 636.990 500.070 637.860 500.210 ;
        RECT 636.990 500.000 637.270 500.070 ;
        RECT 637.720 448.570 637.860 500.070 ;
        RECT 637.260 448.430 637.860 448.570 ;
        RECT 637.260 99.950 637.400 448.430 ;
        RECT 637.200 99.630 637.460 99.950 ;
        RECT 2808.400 99.630 2808.660 99.950 ;
        RECT 2808.460 82.870 2808.600 99.630 ;
        RECT 2808.460 82.730 2809.520 82.870 ;
        RECT 2809.380 2.400 2809.520 82.730 ;
        RECT 2809.170 -4.800 2809.730 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.470 183.500 478.790 183.560 ;
        RECT 904.430 183.500 904.750 183.560 ;
        RECT 478.470 183.360 904.750 183.500 ;
        RECT 478.470 183.300 478.790 183.360 ;
        RECT 904.430 183.300 904.750 183.360 ;
      LAYER via ;
        RECT 478.500 183.300 478.760 183.560 ;
        RECT 904.460 183.300 904.720 183.560 ;
      LAYER met2 ;
        RECT 478.290 500.000 478.570 504.000 ;
        RECT 478.330 499.815 478.470 500.000 ;
        RECT 478.260 499.445 478.540 499.815 ;
        RECT 478.260 498.680 478.540 498.965 ;
        RECT 478.260 498.595 478.700 498.680 ;
        RECT 478.330 498.540 478.700 498.595 ;
        RECT 478.560 183.590 478.700 498.540 ;
        RECT 478.500 183.270 478.760 183.590 ;
        RECT 904.460 183.270 904.720 183.590 ;
        RECT 904.520 82.870 904.660 183.270 ;
        RECT 904.520 82.730 905.120 82.870 ;
        RECT 904.980 2.400 905.120 82.730 ;
        RECT 904.770 -4.800 905.330 2.400 ;
      LAYER via2 ;
        RECT 478.260 499.490 478.540 499.770 ;
        RECT 478.260 498.640 478.540 498.920 ;
      LAYER met3 ;
        RECT 478.235 499.780 478.565 499.795 ;
        RECT 478.020 499.465 478.565 499.780 ;
        RECT 478.020 498.945 478.320 499.465 ;
        RECT 478.020 498.630 478.565 498.945 ;
        RECT 478.235 498.615 478.565 498.630 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 479.620 499.500 479.940 499.760 ;
        RECT 479.710 499.360 479.850 499.500 ;
        RECT 479.480 499.220 479.850 499.360 ;
        RECT 479.480 498.400 479.620 499.220 ;
        RECT 479.390 498.140 479.710 498.400 ;
        RECT 479.390 473.520 479.710 473.580 ;
        RECT 481.690 473.520 482.010 473.580 ;
        RECT 479.390 473.380 482.010 473.520 ;
        RECT 479.390 473.320 479.710 473.380 ;
        RECT 481.690 473.320 482.010 473.380 ;
        RECT 481.690 94.420 482.010 94.480 ;
        RECT 917.770 94.420 918.090 94.480 ;
        RECT 481.690 94.280 918.090 94.420 ;
        RECT 481.690 94.220 482.010 94.280 ;
        RECT 917.770 94.220 918.090 94.280 ;
      LAYER via ;
        RECT 479.650 499.500 479.910 499.760 ;
        RECT 479.420 498.140 479.680 498.400 ;
        RECT 479.420 473.320 479.680 473.580 ;
        RECT 481.720 473.320 481.980 473.580 ;
        RECT 481.720 94.220 481.980 94.480 ;
        RECT 917.800 94.220 918.060 94.480 ;
      LAYER met2 ;
        RECT 479.670 500.000 479.950 504.000 ;
        RECT 479.710 499.790 479.850 500.000 ;
        RECT 479.650 499.470 479.910 499.790 ;
        RECT 479.420 498.110 479.680 498.430 ;
        RECT 479.480 473.610 479.620 498.110 ;
        RECT 479.420 473.290 479.680 473.610 ;
        RECT 481.720 473.290 481.980 473.610 ;
        RECT 481.780 94.510 481.920 473.290 ;
        RECT 481.720 94.190 481.980 94.510 ;
        RECT 917.800 94.190 918.060 94.510 ;
        RECT 917.860 82.870 918.000 94.190 ;
        RECT 917.860 82.730 921.680 82.870 ;
        RECT 921.540 2.400 921.680 82.730 ;
        RECT 921.330 -4.800 921.890 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 16.900 931.890 16.960 ;
        RECT 938.010 16.900 938.330 16.960 ;
        RECT 931.570 16.760 938.330 16.900 ;
        RECT 931.570 16.700 931.890 16.760 ;
        RECT 938.010 16.700 938.330 16.760 ;
      LAYER via ;
        RECT 931.600 16.700 931.860 16.960 ;
        RECT 938.040 16.700 938.300 16.960 ;
      LAYER met2 ;
        RECT 481.050 500.000 481.330 504.000 ;
        RECT 481.090 499.645 481.230 500.000 ;
        RECT 481.020 499.275 481.300 499.645 ;
        RECT 931.590 185.795 931.870 186.165 ;
        RECT 931.660 16.990 931.800 185.795 ;
        RECT 931.600 16.670 931.860 16.990 ;
        RECT 938.040 16.670 938.300 16.990 ;
        RECT 938.100 2.400 938.240 16.670 ;
        RECT 937.890 -4.800 938.450 2.400 ;
      LAYER via2 ;
        RECT 481.020 499.320 481.300 499.600 ;
        RECT 931.590 185.840 931.870 186.120 ;
      LAYER met3 ;
        RECT 479.590 499.610 479.970 499.620 ;
        RECT 480.995 499.610 481.325 499.625 ;
        RECT 479.590 499.310 481.325 499.610 ;
        RECT 479.590 499.300 479.970 499.310 ;
        RECT 480.995 499.295 481.325 499.310 ;
        RECT 479.590 186.130 479.970 186.140 ;
        RECT 931.565 186.130 931.895 186.145 ;
        RECT 479.590 185.830 931.895 186.130 ;
        RECT 479.590 185.820 479.970 185.830 ;
        RECT 931.565 185.815 931.895 185.830 ;
      LAYER via3 ;
        RECT 479.620 499.300 479.940 499.620 ;
        RECT 479.620 185.820 479.940 186.140 ;
      LAYER met4 ;
        RECT 479.615 499.295 479.945 499.625 ;
        RECT 479.630 186.145 479.930 499.295 ;
        RECT 479.615 185.815 479.945 186.145 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.430 500.000 482.710 504.000 ;
        RECT 482.470 498.340 482.610 500.000 ;
        RECT 482.470 498.200 482.840 498.340 ;
        RECT 482.700 488.085 482.840 498.200 ;
        RECT 482.630 487.715 482.910 488.085 ;
        RECT 952.290 202.795 952.570 203.165 ;
        RECT 952.360 82.870 952.500 202.795 ;
        RECT 952.360 82.730 954.800 82.870 ;
        RECT 954.660 2.400 954.800 82.730 ;
        RECT 954.450 -4.800 955.010 2.400 ;
      LAYER via2 ;
        RECT 482.630 487.760 482.910 488.040 ;
        RECT 952.290 202.840 952.570 203.120 ;
      LAYER met3 ;
        RECT 478.670 488.050 479.050 488.060 ;
        RECT 482.605 488.050 482.935 488.065 ;
        RECT 478.670 487.750 482.935 488.050 ;
        RECT 478.670 487.740 479.050 487.750 ;
        RECT 482.605 487.735 482.935 487.750 ;
        RECT 478.670 203.130 479.050 203.140 ;
        RECT 952.265 203.130 952.595 203.145 ;
        RECT 478.670 202.830 952.595 203.130 ;
        RECT 478.670 202.820 479.050 202.830 ;
        RECT 952.265 202.815 952.595 202.830 ;
      LAYER via3 ;
        RECT 478.700 487.740 479.020 488.060 ;
        RECT 478.700 202.820 479.020 203.140 ;
      LAYER met4 ;
        RECT 478.695 487.735 479.025 488.065 ;
        RECT 478.710 203.145 479.010 487.735 ;
        RECT 478.695 202.815 479.025 203.145 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 481.340 483.390 481.400 ;
        RECT 966.070 481.340 966.390 481.400 ;
        RECT 483.070 481.200 966.390 481.340 ;
        RECT 483.070 481.140 483.390 481.200 ;
        RECT 966.070 481.140 966.390 481.200 ;
      LAYER via ;
        RECT 483.100 481.140 483.360 481.400 ;
        RECT 966.100 481.140 966.360 481.400 ;
      LAYER met2 ;
        RECT 483.810 500.000 484.090 504.000 ;
        RECT 483.850 499.645 483.990 500.000 ;
        RECT 483.780 499.275 484.060 499.645 ;
        RECT 483.090 497.915 483.370 498.285 ;
        RECT 483.160 481.430 483.300 497.915 ;
        RECT 483.100 481.110 483.360 481.430 ;
        RECT 966.100 481.110 966.360 481.430 ;
        RECT 966.160 82.870 966.300 481.110 ;
        RECT 966.160 82.730 971.360 82.870 ;
        RECT 971.220 2.400 971.360 82.730 ;
        RECT 971.010 -4.800 971.570 2.400 ;
      LAYER via2 ;
        RECT 483.780 499.320 484.060 499.600 ;
        RECT 483.090 497.960 483.370 498.240 ;
      LAYER met3 ;
        RECT 483.755 499.610 484.085 499.625 ;
        RECT 482.850 499.310 484.085 499.610 ;
        RECT 482.850 498.265 483.150 499.310 ;
        RECT 483.755 499.295 484.085 499.310 ;
        RECT 482.850 497.950 483.395 498.265 ;
        RECT 483.065 497.935 483.395 497.950 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.910 183.160 485.230 183.220 ;
        RECT 987.230 183.160 987.550 183.220 ;
        RECT 484.910 183.020 987.550 183.160 ;
        RECT 484.910 182.960 485.230 183.020 ;
        RECT 987.230 182.960 987.550 183.020 ;
      LAYER via ;
        RECT 484.940 182.960 485.200 183.220 ;
        RECT 987.260 182.960 987.520 183.220 ;
      LAYER met2 ;
        RECT 485.190 500.000 485.470 504.000 ;
        RECT 485.230 499.815 485.370 500.000 ;
        RECT 485.160 499.445 485.440 499.815 ;
        RECT 484.930 497.915 485.210 498.285 ;
        RECT 485.000 183.250 485.140 497.915 ;
        RECT 484.940 182.930 485.200 183.250 ;
        RECT 987.260 182.930 987.520 183.250 ;
        RECT 987.320 82.870 987.460 182.930 ;
        RECT 987.320 82.730 987.920 82.870 ;
        RECT 987.780 2.400 987.920 82.730 ;
        RECT 987.570 -4.800 988.130 2.400 ;
      LAYER via2 ;
        RECT 485.160 499.490 485.440 499.770 ;
        RECT 484.930 497.960 485.210 498.240 ;
      LAYER met3 ;
        RECT 485.135 499.465 485.465 499.795 ;
        RECT 485.150 498.265 485.450 499.465 ;
        RECT 484.905 497.950 485.450 498.265 ;
        RECT 484.905 497.935 485.235 497.950 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 486.520 499.160 486.840 499.420 ;
        RECT 486.610 498.000 486.750 499.160 ;
        RECT 487.210 498.000 487.530 498.060 ;
        RECT 486.610 497.860 487.530 498.000 ;
        RECT 487.210 497.800 487.530 497.860 ;
        RECT 487.210 481.000 487.530 481.060 ;
        RECT 1000.570 481.000 1000.890 481.060 ;
        RECT 487.210 480.860 1000.890 481.000 ;
        RECT 487.210 480.800 487.530 480.860 ;
        RECT 1000.570 480.800 1000.890 480.860 ;
      LAYER via ;
        RECT 486.550 499.160 486.810 499.420 ;
        RECT 487.240 497.800 487.500 498.060 ;
        RECT 487.240 480.800 487.500 481.060 ;
        RECT 1000.600 480.800 1000.860 481.060 ;
      LAYER met2 ;
        RECT 486.570 500.000 486.850 504.000 ;
        RECT 486.610 499.450 486.750 500.000 ;
        RECT 486.550 499.130 486.810 499.450 ;
        RECT 487.240 497.770 487.500 498.090 ;
        RECT 487.300 481.090 487.440 497.770 ;
        RECT 487.240 480.770 487.500 481.090 ;
        RECT 1000.600 480.770 1000.860 481.090 ;
        RECT 1000.660 82.870 1000.800 480.770 ;
        RECT 1000.660 82.730 1004.480 82.870 ;
        RECT 1004.340 2.400 1004.480 82.730 ;
        RECT 1004.130 -4.800 1004.690 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.900 500.860 488.220 501.120 ;
        RECT 487.990 498.400 488.130 500.860 ;
        RECT 487.990 498.200 488.450 498.400 ;
        RECT 488.130 498.140 488.450 498.200 ;
        RECT 1014.370 16.900 1014.690 16.960 ;
        RECT 1020.810 16.900 1021.130 16.960 ;
        RECT 1014.370 16.760 1021.130 16.900 ;
        RECT 1014.370 16.700 1014.690 16.760 ;
        RECT 1020.810 16.700 1021.130 16.760 ;
      LAYER via ;
        RECT 487.930 500.860 488.190 501.120 ;
        RECT 488.160 498.140 488.420 498.400 ;
        RECT 1014.400 16.700 1014.660 16.960 ;
        RECT 1020.840 16.700 1021.100 16.960 ;
      LAYER met2 ;
        RECT 487.950 501.150 488.230 504.000 ;
        RECT 487.930 500.830 488.230 501.150 ;
        RECT 487.950 500.000 488.230 500.830 ;
        RECT 488.160 498.110 488.420 498.430 ;
        RECT 488.220 487.405 488.360 498.110 ;
        RECT 488.150 487.035 488.430 487.405 ;
        RECT 1014.390 185.115 1014.670 185.485 ;
        RECT 1014.460 16.990 1014.600 185.115 ;
        RECT 1014.400 16.670 1014.660 16.990 ;
        RECT 1020.840 16.670 1021.100 16.990 ;
        RECT 1020.900 2.400 1021.040 16.670 ;
        RECT 1020.690 -4.800 1021.250 2.400 ;
      LAYER via2 ;
        RECT 488.150 487.080 488.430 487.360 ;
        RECT 1014.390 185.160 1014.670 185.440 ;
      LAYER met3 ;
        RECT 486.950 487.370 487.330 487.380 ;
        RECT 488.125 487.370 488.455 487.385 ;
        RECT 486.950 487.070 488.455 487.370 ;
        RECT 486.950 487.060 487.330 487.070 ;
        RECT 488.125 487.055 488.455 487.070 ;
        RECT 486.950 185.450 487.330 185.460 ;
        RECT 1014.365 185.450 1014.695 185.465 ;
        RECT 486.950 185.150 1014.695 185.450 ;
        RECT 486.950 185.140 487.330 185.150 ;
        RECT 1014.365 185.135 1014.695 185.150 ;
      LAYER via3 ;
        RECT 486.980 487.060 487.300 487.380 ;
        RECT 486.980 185.140 487.300 185.460 ;
      LAYER met4 ;
        RECT 486.975 487.055 487.305 487.385 ;
        RECT 486.990 185.465 487.290 487.055 ;
        RECT 486.975 185.135 487.305 185.465 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.830 471.820 463.150 471.880 ;
        RECT 465.130 471.820 465.450 471.880 ;
        RECT 462.830 471.680 465.450 471.820 ;
        RECT 462.830 471.620 463.150 471.680 ;
        RECT 465.130 471.620 465.450 471.680 ;
        RECT 465.130 88.300 465.450 88.360 ;
        RECT 717.670 88.300 717.990 88.360 ;
        RECT 465.130 88.160 717.990 88.300 ;
        RECT 465.130 88.100 465.450 88.160 ;
        RECT 717.670 88.100 717.990 88.160 ;
      LAYER via ;
        RECT 462.860 471.620 463.120 471.880 ;
        RECT 465.160 471.620 465.420 471.880 ;
        RECT 465.160 88.100 465.420 88.360 ;
        RECT 717.700 88.100 717.960 88.360 ;
      LAYER met2 ;
        RECT 463.110 500.000 463.390 504.000 ;
        RECT 463.150 499.815 463.290 500.000 ;
        RECT 463.080 499.445 463.360 499.815 ;
        RECT 462.850 497.915 463.130 498.285 ;
        RECT 462.920 471.910 463.060 497.915 ;
        RECT 462.860 471.590 463.120 471.910 ;
        RECT 465.160 471.590 465.420 471.910 ;
        RECT 465.220 88.390 465.360 471.590 ;
        RECT 465.160 88.070 465.420 88.390 ;
        RECT 717.700 88.070 717.960 88.390 ;
        RECT 717.760 82.870 717.900 88.070 ;
        RECT 717.760 82.730 722.960 82.870 ;
        RECT 722.820 2.400 722.960 82.730 ;
        RECT 722.610 -4.800 723.170 2.400 ;
      LAYER via2 ;
        RECT 463.080 499.490 463.360 499.770 ;
        RECT 462.850 497.960 463.130 498.240 ;
      LAYER met3 ;
        RECT 463.055 499.465 463.385 499.795 ;
        RECT 463.070 498.265 463.370 499.465 ;
        RECT 462.825 497.950 463.370 498.265 ;
        RECT 462.825 497.935 463.155 497.950 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.330 500.000 489.610 504.000 ;
        RECT 489.370 498.680 489.510 500.000 ;
        RECT 489.140 498.540 489.510 498.680 ;
        RECT 489.140 486.045 489.280 498.540 ;
        RECT 489.070 485.675 489.350 486.045 ;
        RECT 1035.090 191.235 1035.370 191.605 ;
        RECT 1035.160 82.870 1035.300 191.235 ;
        RECT 1035.160 82.730 1037.600 82.870 ;
        RECT 1037.460 2.400 1037.600 82.730 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
      LAYER via2 ;
        RECT 489.070 485.720 489.350 486.000 ;
        RECT 1035.090 191.280 1035.370 191.560 ;
      LAYER met3 ;
        RECT 486.030 486.010 486.410 486.020 ;
        RECT 489.045 486.010 489.375 486.025 ;
        RECT 486.030 485.710 489.375 486.010 ;
        RECT 486.030 485.700 486.410 485.710 ;
        RECT 489.045 485.695 489.375 485.710 ;
        RECT 486.030 191.570 486.410 191.580 ;
        RECT 1035.065 191.570 1035.395 191.585 ;
        RECT 486.030 191.270 1035.395 191.570 ;
        RECT 486.030 191.260 486.410 191.270 ;
        RECT 1035.065 191.255 1035.395 191.270 ;
      LAYER via3 ;
        RECT 486.060 485.700 486.380 486.020 ;
        RECT 486.060 191.260 486.380 191.580 ;
      LAYER met4 ;
        RECT 486.055 485.695 486.385 486.025 ;
        RECT 486.070 191.585 486.370 485.695 ;
        RECT 486.055 191.255 486.385 191.585 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.660 498.820 490.980 499.080 ;
        RECT 490.750 496.980 490.890 498.820 ;
        RECT 505.150 496.980 505.470 497.040 ;
        RECT 490.750 496.840 505.470 496.980 ;
        RECT 505.150 496.780 505.470 496.840 ;
        RECT 505.150 482.020 505.470 482.080 ;
        RECT 679.950 482.020 680.270 482.080 ;
        RECT 505.150 481.880 680.270 482.020 ;
        RECT 505.150 481.820 505.470 481.880 ;
        RECT 679.950 481.820 680.270 481.880 ;
        RECT 807.230 19.820 821.860 19.960 ;
        RECT 679.950 19.620 680.270 19.680 ;
        RECT 807.230 19.620 807.370 19.820 ;
        RECT 679.950 19.480 807.370 19.620 ;
        RECT 821.720 19.620 821.860 19.820 ;
        RECT 1053.930 19.620 1054.250 19.680 ;
        RECT 821.720 19.480 1054.250 19.620 ;
        RECT 679.950 19.420 680.270 19.480 ;
        RECT 1053.930 19.420 1054.250 19.480 ;
      LAYER via ;
        RECT 490.690 498.820 490.950 499.080 ;
        RECT 505.180 496.780 505.440 497.040 ;
        RECT 505.180 481.820 505.440 482.080 ;
        RECT 679.980 481.820 680.240 482.080 ;
        RECT 679.980 19.420 680.240 19.680 ;
        RECT 1053.960 19.420 1054.220 19.680 ;
      LAYER met2 ;
        RECT 490.710 500.000 490.990 504.000 ;
        RECT 490.750 499.110 490.890 500.000 ;
        RECT 490.690 498.790 490.950 499.110 ;
        RECT 505.180 496.750 505.440 497.070 ;
        RECT 505.240 482.110 505.380 496.750 ;
        RECT 505.180 481.790 505.440 482.110 ;
        RECT 679.980 481.790 680.240 482.110 ;
        RECT 680.040 19.710 680.180 481.790 ;
        RECT 679.980 19.390 680.240 19.710 ;
        RECT 1053.960 19.390 1054.220 19.710 ;
        RECT 1054.020 2.400 1054.160 19.390 ;
        RECT 1053.810 -4.800 1054.370 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.040 499.700 492.360 499.760 ;
        RECT 491.900 499.500 492.360 499.700 ;
        RECT 491.900 498.740 492.040 499.500 ;
        RECT 491.810 498.480 492.130 498.740 ;
        RECT 489.970 473.180 490.290 473.240 ;
        RECT 491.810 473.180 492.130 473.240 ;
        RECT 489.970 473.040 492.130 473.180 ;
        RECT 489.970 472.980 490.290 473.040 ;
        RECT 491.810 472.980 492.130 473.040 ;
        RECT 489.970 102.240 490.290 102.300 ;
        RECT 1069.570 102.240 1069.890 102.300 ;
        RECT 489.970 102.100 1069.890 102.240 ;
        RECT 489.970 102.040 490.290 102.100 ;
        RECT 1069.570 102.040 1069.890 102.100 ;
      LAYER via ;
        RECT 492.070 499.500 492.330 499.760 ;
        RECT 491.840 498.480 492.100 498.740 ;
        RECT 490.000 472.980 490.260 473.240 ;
        RECT 491.840 472.980 492.100 473.240 ;
        RECT 490.000 102.040 490.260 102.300 ;
        RECT 1069.600 102.040 1069.860 102.300 ;
      LAYER met2 ;
        RECT 492.090 500.000 492.370 504.000 ;
        RECT 492.130 499.790 492.270 500.000 ;
        RECT 492.070 499.470 492.330 499.790 ;
        RECT 491.840 498.450 492.100 498.770 ;
        RECT 491.900 473.270 492.040 498.450 ;
        RECT 490.000 472.950 490.260 473.270 ;
        RECT 491.840 472.950 492.100 473.270 ;
        RECT 490.060 102.330 490.200 472.950 ;
        RECT 490.000 102.010 490.260 102.330 ;
        RECT 1069.600 102.010 1069.860 102.330 ;
        RECT 1069.660 82.870 1069.800 102.010 ;
        RECT 1069.660 82.730 1070.720 82.870 ;
        RECT 1070.580 2.400 1070.720 82.730 ;
        RECT 1070.370 -4.800 1070.930 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 493.420 499.500 493.740 499.760 ;
        RECT 493.510 498.740 493.650 499.500 ;
        RECT 493.510 498.540 493.970 498.740 ;
        RECT 493.650 498.480 493.970 498.540 ;
        RECT 491.810 471.820 492.130 471.880 ;
        RECT 493.650 471.820 493.970 471.880 ;
        RECT 491.810 471.680 493.970 471.820 ;
        RECT 491.810 471.620 492.130 471.680 ;
        RECT 493.650 471.620 493.970 471.680 ;
        RECT 491.810 164.460 492.130 164.520 ;
        RECT 1083.370 164.460 1083.690 164.520 ;
        RECT 491.810 164.320 1083.690 164.460 ;
        RECT 491.810 164.260 492.130 164.320 ;
        RECT 1083.370 164.260 1083.690 164.320 ;
      LAYER via ;
        RECT 493.450 499.500 493.710 499.760 ;
        RECT 493.680 498.480 493.940 498.740 ;
        RECT 491.840 471.620 492.100 471.880 ;
        RECT 493.680 471.620 493.940 471.880 ;
        RECT 491.840 164.260 492.100 164.520 ;
        RECT 1083.400 164.260 1083.660 164.520 ;
      LAYER met2 ;
        RECT 493.470 500.000 493.750 504.000 ;
        RECT 493.510 499.790 493.650 500.000 ;
        RECT 493.450 499.470 493.710 499.790 ;
        RECT 493.680 498.450 493.940 498.770 ;
        RECT 493.740 471.910 493.880 498.450 ;
        RECT 491.840 471.590 492.100 471.910 ;
        RECT 493.680 471.590 493.940 471.910 ;
        RECT 491.900 164.550 492.040 471.590 ;
        RECT 491.840 164.230 492.100 164.550 ;
        RECT 1083.400 164.230 1083.660 164.550 ;
        RECT 1083.460 82.870 1083.600 164.230 ;
        RECT 1083.460 82.730 1087.280 82.870 ;
        RECT 1087.140 2.400 1087.280 82.730 ;
        RECT 1086.930 -4.800 1087.490 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 494.800 500.720 495.120 500.780 ;
        RECT 493.050 500.580 495.120 500.720 ;
        RECT 493.050 497.320 493.190 500.580 ;
        RECT 494.800 500.520 495.120 500.580 ;
        RECT 495.030 497.320 495.350 497.380 ;
        RECT 493.050 497.180 495.350 497.320 ;
        RECT 495.030 497.120 495.350 497.180 ;
        RECT 1097.630 19.620 1097.950 19.680 ;
        RECT 1103.610 19.620 1103.930 19.680 ;
        RECT 1097.630 19.480 1103.930 19.620 ;
        RECT 1097.630 19.420 1097.950 19.480 ;
        RECT 1103.610 19.420 1103.930 19.480 ;
      LAYER via ;
        RECT 494.830 500.520 495.090 500.780 ;
        RECT 495.060 497.120 495.320 497.380 ;
        RECT 1097.660 19.420 1097.920 19.680 ;
        RECT 1103.640 19.420 1103.900 19.680 ;
      LAYER met2 ;
        RECT 494.850 500.810 495.130 504.000 ;
        RECT 494.830 500.490 495.130 500.810 ;
        RECT 494.850 500.000 495.130 500.490 ;
        RECT 495.060 497.090 495.320 497.410 ;
        RECT 495.120 487.405 495.260 497.090 ;
        RECT 495.050 487.035 495.330 487.405 ;
        RECT 1097.650 106.915 1097.930 107.285 ;
        RECT 1097.720 19.710 1097.860 106.915 ;
        RECT 1097.660 19.390 1097.920 19.710 ;
        RECT 1103.640 19.390 1103.900 19.710 ;
        RECT 1103.700 2.400 1103.840 19.390 ;
        RECT 1103.490 -4.800 1104.050 2.400 ;
      LAYER via2 ;
        RECT 495.050 487.080 495.330 487.360 ;
        RECT 1097.650 106.960 1097.930 107.240 ;
      LAYER met3 ;
        RECT 495.025 487.380 495.355 487.385 ;
        RECT 495.025 487.370 495.610 487.380 ;
        RECT 495.025 487.070 495.810 487.370 ;
        RECT 495.025 487.060 495.610 487.070 ;
        RECT 495.025 487.055 495.355 487.060 ;
        RECT 495.230 107.250 495.610 107.260 ;
        RECT 1097.625 107.250 1097.955 107.265 ;
        RECT 495.230 106.950 1097.955 107.250 ;
        RECT 495.230 106.940 495.610 106.950 ;
        RECT 1097.625 106.935 1097.955 106.950 ;
      LAYER via3 ;
        RECT 495.260 487.060 495.580 487.380 ;
        RECT 495.260 106.940 495.580 107.260 ;
      LAYER met4 ;
        RECT 495.255 487.055 495.585 487.385 ;
        RECT 495.270 107.265 495.570 487.055 ;
        RECT 495.255 106.935 495.585 107.265 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.180 499.160 496.500 499.420 ;
        RECT 494.110 498.000 494.430 498.060 ;
        RECT 496.270 498.000 496.410 499.160 ;
        RECT 494.110 497.860 496.410 498.000 ;
        RECT 494.110 497.800 494.430 497.860 ;
      LAYER via ;
        RECT 496.210 499.160 496.470 499.420 ;
        RECT 494.140 497.800 494.400 498.060 ;
      LAYER met2 ;
        RECT 496.230 500.000 496.510 504.000 ;
        RECT 496.270 499.450 496.410 500.000 ;
        RECT 496.210 499.130 496.470 499.450 ;
        RECT 494.140 497.770 494.400 498.090 ;
        RECT 494.200 497.605 494.340 497.770 ;
        RECT 494.130 497.235 494.410 497.605 ;
        RECT 1117.890 190.555 1118.170 190.925 ;
        RECT 1117.960 82.870 1118.100 190.555 ;
        RECT 1117.960 82.730 1120.400 82.870 ;
        RECT 1120.260 2.400 1120.400 82.730 ;
        RECT 1120.050 -4.800 1120.610 2.400 ;
      LAYER via2 ;
        RECT 494.130 497.280 494.410 497.560 ;
        RECT 1117.890 190.600 1118.170 190.880 ;
      LAYER met3 ;
        RECT 493.390 497.570 493.770 497.580 ;
        RECT 494.105 497.570 494.435 497.585 ;
        RECT 493.390 497.270 494.435 497.570 ;
        RECT 493.390 497.260 493.770 497.270 ;
        RECT 494.105 497.255 494.435 497.270 ;
        RECT 493.390 190.890 493.770 190.900 ;
        RECT 1117.865 190.890 1118.195 190.905 ;
        RECT 493.390 190.590 1118.195 190.890 ;
        RECT 493.390 190.580 493.770 190.590 ;
        RECT 1117.865 190.575 1118.195 190.590 ;
      LAYER via3 ;
        RECT 493.420 497.260 493.740 497.580 ;
        RECT 493.420 190.580 493.740 190.900 ;
      LAYER met4 ;
        RECT 493.415 497.255 493.745 497.585 ;
        RECT 493.430 190.905 493.730 497.255 ;
        RECT 493.415 190.575 493.745 190.905 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.560 499.500 497.880 499.760 ;
        RECT 497.650 498.740 497.790 499.500 ;
        RECT 497.650 498.540 498.110 498.740 ;
        RECT 497.790 498.480 498.110 498.540 ;
        RECT 497.790 108.700 498.110 108.760 ;
        RECT 1131.670 108.700 1131.990 108.760 ;
        RECT 497.790 108.560 1131.990 108.700 ;
        RECT 497.790 108.500 498.110 108.560 ;
        RECT 1131.670 108.500 1131.990 108.560 ;
      LAYER via ;
        RECT 497.590 499.500 497.850 499.760 ;
        RECT 497.820 498.480 498.080 498.740 ;
        RECT 497.820 108.500 498.080 108.760 ;
        RECT 1131.700 108.500 1131.960 108.760 ;
      LAYER met2 ;
        RECT 497.610 500.000 497.890 504.000 ;
        RECT 497.650 499.790 497.790 500.000 ;
        RECT 497.590 499.470 497.850 499.790 ;
        RECT 497.820 498.450 498.080 498.770 ;
        RECT 497.880 108.790 498.020 498.450 ;
        RECT 497.820 108.470 498.080 108.790 ;
        RECT 1131.700 108.470 1131.960 108.790 ;
        RECT 1131.760 82.870 1131.900 108.470 ;
        RECT 1131.760 82.730 1136.960 82.870 ;
        RECT 1136.820 2.400 1136.960 82.730 ;
        RECT 1136.610 -4.800 1137.170 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.250 191.320 498.570 191.380 ;
        RECT 1152.370 191.320 1152.690 191.380 ;
        RECT 498.250 191.180 1152.690 191.320 ;
        RECT 498.250 191.120 498.570 191.180 ;
        RECT 1152.370 191.120 1152.690 191.180 ;
      LAYER via ;
        RECT 498.280 191.120 498.540 191.380 ;
        RECT 1152.400 191.120 1152.660 191.380 ;
      LAYER met2 ;
        RECT 498.990 500.000 499.270 504.000 ;
        RECT 499.030 498.340 499.170 500.000 ;
        RECT 498.340 498.200 499.170 498.340 ;
        RECT 498.340 191.410 498.480 498.200 ;
        RECT 498.280 191.090 498.540 191.410 ;
        RECT 1152.400 191.090 1152.660 191.410 ;
        RECT 1152.460 82.870 1152.600 191.090 ;
        RECT 1152.460 82.730 1153.520 82.870 ;
        RECT 1153.380 2.400 1153.520 82.730 ;
        RECT 1153.170 -4.800 1153.730 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.320 499.160 500.640 499.420 ;
        RECT 500.410 498.680 500.550 499.160 ;
        RECT 500.410 498.540 500.780 498.680 ;
        RECT 498.710 497.660 499.030 497.720 ;
        RECT 500.640 497.660 500.780 498.540 ;
        RECT 498.710 497.520 500.780 497.660 ;
        RECT 498.710 497.460 499.030 497.520 ;
        RECT 498.710 190.980 499.030 191.040 ;
        RECT 1166.170 190.980 1166.490 191.040 ;
        RECT 498.710 190.840 1166.490 190.980 ;
        RECT 498.710 190.780 499.030 190.840 ;
        RECT 1166.170 190.780 1166.490 190.840 ;
      LAYER via ;
        RECT 500.350 499.160 500.610 499.420 ;
        RECT 498.740 497.460 499.000 497.720 ;
        RECT 498.740 190.780 499.000 191.040 ;
        RECT 1166.200 190.780 1166.460 191.040 ;
      LAYER met2 ;
        RECT 500.370 500.000 500.650 504.000 ;
        RECT 500.410 499.450 500.550 500.000 ;
        RECT 500.350 499.130 500.610 499.450 ;
        RECT 498.740 497.430 499.000 497.750 ;
        RECT 498.800 191.070 498.940 497.430 ;
        RECT 498.740 190.750 499.000 191.070 ;
        RECT 1166.200 190.750 1166.460 191.070 ;
        RECT 1166.260 82.870 1166.400 190.750 ;
        RECT 1166.260 82.730 1170.080 82.870 ;
        RECT 1169.940 2.400 1170.080 82.730 ;
        RECT 1169.730 -4.800 1170.290 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1179.970 16.900 1180.290 16.960 ;
        RECT 1186.410 16.900 1186.730 16.960 ;
        RECT 1179.970 16.760 1186.730 16.900 ;
        RECT 1179.970 16.700 1180.290 16.760 ;
        RECT 1186.410 16.700 1186.730 16.760 ;
      LAYER via ;
        RECT 1180.000 16.700 1180.260 16.960 ;
        RECT 1186.440 16.700 1186.700 16.960 ;
      LAYER met2 ;
        RECT 501.750 500.000 502.030 504.000 ;
        RECT 501.790 499.645 501.930 500.000 ;
        RECT 501.720 499.275 502.000 499.645 ;
        RECT 1179.990 472.755 1180.270 473.125 ;
        RECT 1180.060 16.990 1180.200 472.755 ;
        RECT 1180.000 16.670 1180.260 16.990 ;
        RECT 1186.440 16.670 1186.700 16.990 ;
        RECT 1186.500 2.400 1186.640 16.670 ;
        RECT 1186.290 -4.800 1186.850 2.400 ;
      LAYER via2 ;
        RECT 501.720 499.320 502.000 499.600 ;
        RECT 1179.990 472.800 1180.270 473.080 ;
      LAYER met3 ;
        RECT 501.695 499.610 502.025 499.625 ;
        RECT 502.590 499.610 502.970 499.620 ;
        RECT 501.695 499.310 502.970 499.610 ;
        RECT 501.695 499.295 502.025 499.310 ;
        RECT 502.590 499.300 502.970 499.310 ;
        RECT 502.590 473.090 502.970 473.100 ;
        RECT 1179.965 473.090 1180.295 473.105 ;
        RECT 502.590 472.790 1180.295 473.090 ;
        RECT 502.590 472.780 502.970 472.790 ;
        RECT 1179.965 472.775 1180.295 472.790 ;
      LAYER via3 ;
        RECT 502.620 499.300 502.940 499.620 ;
        RECT 502.620 472.780 502.940 473.100 ;
      LAYER met4 ;
        RECT 502.615 499.295 502.945 499.625 ;
        RECT 502.630 473.105 502.930 499.295 ;
        RECT 502.615 472.775 502.945 473.105 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.440 499.500 464.760 499.760 ;
        RECT 464.530 498.740 464.670 499.500 ;
        RECT 464.210 498.540 464.670 498.740 ;
        RECT 464.210 498.480 464.530 498.540 ;
        RECT 464.210 487.800 464.530 487.860 ;
        RECT 467.430 487.800 467.750 487.860 ;
        RECT 464.210 487.660 467.750 487.800 ;
        RECT 464.210 487.600 464.530 487.660 ;
        RECT 467.430 487.600 467.750 487.660 ;
        RECT 467.890 109.380 468.210 109.440 ;
        RECT 738.370 109.380 738.690 109.440 ;
        RECT 467.890 109.240 738.690 109.380 ;
        RECT 467.890 109.180 468.210 109.240 ;
        RECT 738.370 109.180 738.690 109.240 ;
      LAYER via ;
        RECT 464.470 499.500 464.730 499.760 ;
        RECT 464.240 498.480 464.500 498.740 ;
        RECT 464.240 487.600 464.500 487.860 ;
        RECT 467.460 487.600 467.720 487.860 ;
        RECT 467.920 109.180 468.180 109.440 ;
        RECT 738.400 109.180 738.660 109.440 ;
      LAYER met2 ;
        RECT 464.490 500.000 464.770 504.000 ;
        RECT 464.530 499.790 464.670 500.000 ;
        RECT 464.470 499.470 464.730 499.790 ;
        RECT 464.240 498.450 464.500 498.770 ;
        RECT 464.300 487.890 464.440 498.450 ;
        RECT 464.240 487.570 464.500 487.890 ;
        RECT 467.460 487.570 467.720 487.890 ;
        RECT 467.520 448.570 467.660 487.570 ;
        RECT 467.520 448.430 468.120 448.570 ;
        RECT 467.980 109.470 468.120 448.430 ;
        RECT 467.920 109.150 468.180 109.470 ;
        RECT 738.400 109.150 738.660 109.470 ;
        RECT 738.460 17.410 738.600 109.150 ;
        RECT 738.460 17.270 739.520 17.410 ;
        RECT 739.380 2.400 739.520 17.270 ;
        RECT 739.170 -4.800 739.730 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.080 499.500 503.400 499.760 ;
        RECT 503.170 499.080 503.310 499.500 ;
        RECT 503.170 498.880 503.630 499.080 ;
        RECT 503.310 498.820 503.630 498.880 ;
      LAYER via ;
        RECT 503.110 499.500 503.370 499.760 ;
        RECT 503.340 498.820 503.600 499.080 ;
      LAYER met2 ;
        RECT 503.130 500.000 503.410 504.000 ;
        RECT 503.170 499.790 503.310 500.000 ;
        RECT 503.110 499.470 503.370 499.790 ;
        RECT 503.340 498.790 503.600 499.110 ;
        RECT 503.400 492.165 503.540 498.790 ;
        RECT 503.330 491.795 503.610 492.165 ;
        RECT 1200.690 135.475 1200.970 135.845 ;
        RECT 1200.760 82.870 1200.900 135.475 ;
        RECT 1200.760 82.730 1203.200 82.870 ;
        RECT 1203.060 2.400 1203.200 82.730 ;
        RECT 1202.850 -4.800 1203.410 2.400 ;
      LAYER via2 ;
        RECT 503.330 491.840 503.610 492.120 ;
        RECT 1200.690 135.520 1200.970 135.800 ;
      LAYER met3 ;
        RECT 500.750 492.130 501.130 492.140 ;
        RECT 503.305 492.130 503.635 492.145 ;
        RECT 500.750 491.830 503.635 492.130 ;
        RECT 500.750 491.820 501.130 491.830 ;
        RECT 503.305 491.815 503.635 491.830 ;
        RECT 500.750 135.810 501.130 135.820 ;
        RECT 1200.665 135.810 1200.995 135.825 ;
        RECT 500.750 135.510 1200.995 135.810 ;
        RECT 500.750 135.500 501.130 135.510 ;
        RECT 1200.665 135.495 1200.995 135.510 ;
      LAYER via3 ;
        RECT 500.780 491.820 501.100 492.140 ;
        RECT 500.780 135.500 501.100 135.820 ;
      LAYER met4 ;
        RECT 500.775 491.815 501.105 492.145 ;
        RECT 500.790 135.825 501.090 491.815 ;
        RECT 500.775 135.495 501.105 135.825 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.460 499.500 504.780 499.760 ;
        RECT 504.550 498.400 504.690 499.500 ;
        RECT 504.550 498.200 505.010 498.400 ;
        RECT 504.690 498.140 505.010 498.200 ;
        RECT 505.150 472.160 505.470 472.220 ;
        RECT 506.070 472.160 506.390 472.220 ;
        RECT 505.150 472.020 506.390 472.160 ;
        RECT 505.150 471.960 505.470 472.020 ;
        RECT 506.070 471.960 506.390 472.020 ;
        RECT 506.070 205.600 506.390 205.660 ;
        RECT 1214.470 205.600 1214.790 205.660 ;
        RECT 506.070 205.460 1214.790 205.600 ;
        RECT 506.070 205.400 506.390 205.460 ;
        RECT 1214.470 205.400 1214.790 205.460 ;
      LAYER via ;
        RECT 504.490 499.500 504.750 499.760 ;
        RECT 504.720 498.140 504.980 498.400 ;
        RECT 505.180 471.960 505.440 472.220 ;
        RECT 506.100 471.960 506.360 472.220 ;
        RECT 506.100 205.400 506.360 205.660 ;
        RECT 1214.500 205.400 1214.760 205.660 ;
      LAYER met2 ;
        RECT 504.510 500.000 504.790 504.000 ;
        RECT 504.550 499.790 504.690 500.000 ;
        RECT 504.490 499.470 504.750 499.790 ;
        RECT 504.720 498.110 504.980 498.430 ;
        RECT 504.780 473.520 504.920 498.110 ;
        RECT 504.780 473.380 505.380 473.520 ;
        RECT 505.240 472.250 505.380 473.380 ;
        RECT 505.180 471.930 505.440 472.250 ;
        RECT 506.100 471.930 506.360 472.250 ;
        RECT 506.160 205.690 506.300 471.930 ;
        RECT 506.100 205.370 506.360 205.690 ;
        RECT 1214.500 205.370 1214.760 205.690 ;
        RECT 1214.560 82.870 1214.700 205.370 ;
        RECT 1214.560 82.730 1219.760 82.870 ;
        RECT 1219.620 2.400 1219.760 82.730 ;
        RECT 1219.410 -4.800 1219.970 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.070 474.200 506.390 474.260 ;
        RECT 1235.170 474.200 1235.490 474.260 ;
        RECT 506.070 474.060 1235.490 474.200 ;
        RECT 506.070 474.000 506.390 474.060 ;
        RECT 1235.170 474.000 1235.490 474.060 ;
      LAYER via ;
        RECT 506.100 474.000 506.360 474.260 ;
        RECT 1235.200 474.000 1235.460 474.260 ;
      LAYER met2 ;
        RECT 505.890 500.000 506.170 504.000 ;
        RECT 505.930 498.850 506.070 500.000 ;
        RECT 505.930 498.710 506.300 498.850 ;
        RECT 506.160 474.290 506.300 498.710 ;
        RECT 506.100 473.970 506.360 474.290 ;
        RECT 1235.200 473.970 1235.460 474.290 ;
        RECT 1235.260 17.410 1235.400 473.970 ;
        RECT 1235.260 17.270 1236.320 17.410 ;
        RECT 1236.180 2.400 1236.320 17.270 ;
        RECT 1235.970 -4.800 1236.530 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 507.220 499.500 507.540 499.760 ;
        RECT 507.310 499.360 507.450 499.500 ;
        RECT 507.310 499.220 509.060 499.360 ;
        RECT 503.770 497.660 504.090 497.720 ;
        RECT 508.920 497.660 509.060 499.220 ;
        RECT 503.770 497.520 509.060 497.660 ;
        RECT 503.770 497.460 504.090 497.520 ;
        RECT 503.770 114.480 504.090 114.540 ;
        RECT 1248.970 114.480 1249.290 114.540 ;
        RECT 503.770 114.340 1249.290 114.480 ;
        RECT 503.770 114.280 504.090 114.340 ;
        RECT 1248.970 114.280 1249.290 114.340 ;
      LAYER via ;
        RECT 507.250 499.500 507.510 499.760 ;
        RECT 503.800 497.460 504.060 497.720 ;
        RECT 503.800 114.280 504.060 114.540 ;
        RECT 1249.000 114.280 1249.260 114.540 ;
      LAYER met2 ;
        RECT 507.270 500.000 507.550 504.000 ;
        RECT 507.310 499.790 507.450 500.000 ;
        RECT 507.250 499.470 507.510 499.790 ;
        RECT 503.800 497.430 504.060 497.750 ;
        RECT 503.860 114.570 504.000 497.430 ;
        RECT 503.800 114.250 504.060 114.570 ;
        RECT 1249.000 114.250 1249.260 114.570 ;
        RECT 1249.060 82.870 1249.200 114.250 ;
        RECT 1249.060 82.730 1252.880 82.870 ;
        RECT 1252.740 2.400 1252.880 82.730 ;
        RECT 1252.530 -4.800 1253.090 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 508.600 499.700 508.920 499.760 ;
        RECT 508.600 499.560 509.520 499.700 ;
        RECT 508.600 499.500 508.920 499.560 ;
        RECT 509.380 498.060 509.520 499.560 ;
        RECT 509.290 497.800 509.610 498.060 ;
        RECT 509.290 473.860 509.610 473.920 ;
        RECT 1262.770 473.860 1263.090 473.920 ;
        RECT 509.290 473.720 1263.090 473.860 ;
        RECT 509.290 473.660 509.610 473.720 ;
        RECT 1262.770 473.660 1263.090 473.720 ;
        RECT 1262.770 16.900 1263.090 16.960 ;
        RECT 1269.210 16.900 1269.530 16.960 ;
        RECT 1262.770 16.760 1269.530 16.900 ;
        RECT 1262.770 16.700 1263.090 16.760 ;
        RECT 1269.210 16.700 1269.530 16.760 ;
      LAYER via ;
        RECT 508.630 499.500 508.890 499.760 ;
        RECT 509.320 497.800 509.580 498.060 ;
        RECT 509.320 473.660 509.580 473.920 ;
        RECT 1262.800 473.660 1263.060 473.920 ;
        RECT 1262.800 16.700 1263.060 16.960 ;
        RECT 1269.240 16.700 1269.500 16.960 ;
      LAYER met2 ;
        RECT 508.650 500.000 508.930 504.000 ;
        RECT 508.690 499.790 508.830 500.000 ;
        RECT 508.630 499.470 508.890 499.790 ;
        RECT 509.320 497.770 509.580 498.090 ;
        RECT 509.380 473.950 509.520 497.770 ;
        RECT 509.320 473.630 509.580 473.950 ;
        RECT 1262.800 473.630 1263.060 473.950 ;
        RECT 1262.860 16.990 1263.000 473.630 ;
        RECT 1262.800 16.670 1263.060 16.990 ;
        RECT 1269.240 16.670 1269.500 16.990 ;
        RECT 1269.300 2.400 1269.440 16.670 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.030 500.000 510.310 504.000 ;
        RECT 510.070 499.815 510.210 500.000 ;
        RECT 510.000 499.445 510.280 499.815 ;
        RECT 510.230 491.115 510.510 491.485 ;
        RECT 510.300 477.885 510.440 491.115 ;
        RECT 510.230 477.515 510.510 477.885 ;
        RECT 1283.490 114.395 1283.770 114.765 ;
        RECT 1283.560 82.870 1283.700 114.395 ;
        RECT 1283.560 82.730 1286.000 82.870 ;
        RECT 1285.860 2.400 1286.000 82.730 ;
        RECT 1285.650 -4.800 1286.210 2.400 ;
      LAYER via2 ;
        RECT 510.000 499.490 510.280 499.770 ;
        RECT 510.230 491.160 510.510 491.440 ;
        RECT 510.230 477.560 510.510 477.840 ;
        RECT 1283.490 114.440 1283.770 114.720 ;
      LAYER met3 ;
        RECT 509.975 499.610 510.305 499.795 ;
        RECT 510.870 499.610 511.250 499.620 ;
        RECT 509.975 499.465 511.250 499.610 ;
        RECT 509.990 499.310 511.250 499.465 ;
        RECT 510.870 499.300 511.250 499.310 ;
        RECT 510.205 491.450 510.535 491.465 ;
        RECT 510.870 491.450 511.250 491.460 ;
        RECT 510.205 491.150 511.250 491.450 ;
        RECT 510.205 491.135 510.535 491.150 ;
        RECT 510.870 491.140 511.250 491.150 ;
        RECT 509.030 477.850 509.410 477.860 ;
        RECT 510.205 477.850 510.535 477.865 ;
        RECT 509.030 477.550 510.535 477.850 ;
        RECT 509.030 477.540 509.410 477.550 ;
        RECT 510.205 477.535 510.535 477.550 ;
        RECT 509.030 114.730 509.410 114.740 ;
        RECT 1283.465 114.730 1283.795 114.745 ;
        RECT 509.030 114.430 1283.795 114.730 ;
        RECT 509.030 114.420 509.410 114.430 ;
        RECT 1283.465 114.415 1283.795 114.430 ;
      LAYER via3 ;
        RECT 510.900 499.300 511.220 499.620 ;
        RECT 510.900 491.140 511.220 491.460 ;
        RECT 509.060 477.540 509.380 477.860 ;
        RECT 509.060 114.420 509.380 114.740 ;
      LAYER met4 ;
        RECT 510.895 499.295 511.225 499.625 ;
        RECT 510.910 491.465 511.210 499.295 ;
        RECT 510.895 491.135 511.225 491.465 ;
        RECT 509.055 477.535 509.385 477.865 ;
        RECT 509.070 114.745 509.370 477.535 ;
        RECT 509.055 114.415 509.385 114.745 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.360 499.500 511.680 499.760 ;
        RECT 511.450 499.080 511.590 499.500 ;
        RECT 511.450 498.880 511.910 499.080 ;
        RECT 511.590 498.820 511.910 498.880 ;
        RECT 511.130 477.260 511.450 477.320 ;
        RECT 512.970 477.260 513.290 477.320 ;
        RECT 511.130 477.120 513.290 477.260 ;
        RECT 511.130 477.060 511.450 477.120 ;
        RECT 512.970 477.060 513.290 477.120 ;
        RECT 512.970 114.140 513.290 114.200 ;
        RECT 1297.270 114.140 1297.590 114.200 ;
        RECT 512.970 114.000 1297.590 114.140 ;
        RECT 512.970 113.940 513.290 114.000 ;
        RECT 1297.270 113.940 1297.590 114.000 ;
      LAYER via ;
        RECT 511.390 499.500 511.650 499.760 ;
        RECT 511.620 498.820 511.880 499.080 ;
        RECT 511.160 477.060 511.420 477.320 ;
        RECT 513.000 477.060 513.260 477.320 ;
        RECT 513.000 113.940 513.260 114.200 ;
        RECT 1297.300 113.940 1297.560 114.200 ;
      LAYER met2 ;
        RECT 511.410 500.000 511.690 504.000 ;
        RECT 511.450 499.790 511.590 500.000 ;
        RECT 511.390 499.470 511.650 499.790 ;
        RECT 511.620 498.790 511.880 499.110 ;
        RECT 511.680 498.000 511.820 498.790 ;
        RECT 511.220 497.860 511.820 498.000 ;
        RECT 511.220 477.350 511.360 497.860 ;
        RECT 511.160 477.030 511.420 477.350 ;
        RECT 513.000 477.030 513.260 477.350 ;
        RECT 513.060 114.230 513.200 477.030 ;
        RECT 513.000 113.910 513.260 114.230 ;
        RECT 1297.300 113.910 1297.560 114.230 ;
        RECT 1297.360 82.870 1297.500 113.910 ;
        RECT 1297.360 82.730 1302.560 82.870 ;
        RECT 1302.420 2.400 1302.560 82.730 ;
        RECT 1302.210 -4.800 1302.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 512.510 113.800 512.830 113.860 ;
        RECT 1317.970 113.800 1318.290 113.860 ;
        RECT 512.510 113.660 1318.290 113.800 ;
        RECT 512.510 113.600 512.830 113.660 ;
        RECT 1317.970 113.600 1318.290 113.660 ;
      LAYER via ;
        RECT 512.540 113.600 512.800 113.860 ;
        RECT 1318.000 113.600 1318.260 113.860 ;
      LAYER met2 ;
        RECT 512.790 500.000 513.070 504.000 ;
        RECT 512.830 499.815 512.970 500.000 ;
        RECT 512.760 499.445 513.040 499.815 ;
        RECT 512.530 498.595 512.810 498.965 ;
        RECT 512.600 113.890 512.740 498.595 ;
        RECT 512.540 113.570 512.800 113.890 ;
        RECT 1318.000 113.570 1318.260 113.890 ;
        RECT 1318.060 82.870 1318.200 113.570 ;
        RECT 1318.060 82.730 1319.120 82.870 ;
        RECT 1318.980 2.400 1319.120 82.730 ;
        RECT 1318.770 -4.800 1319.330 2.400 ;
      LAYER via2 ;
        RECT 512.760 499.490 513.040 499.770 ;
        RECT 512.530 498.640 512.810 498.920 ;
      LAYER met3 ;
        RECT 512.735 499.465 513.065 499.795 ;
        RECT 512.750 498.945 513.050 499.465 ;
        RECT 512.505 498.630 513.050 498.945 ;
        RECT 512.505 498.615 512.835 498.630 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.120 499.700 514.440 499.760 ;
        RECT 514.120 499.560 515.960 499.700 ;
        RECT 514.120 499.500 514.440 499.560 ;
        RECT 515.820 497.660 515.960 499.560 ;
        RECT 516.650 497.660 516.970 497.720 ;
        RECT 515.820 497.520 516.970 497.660 ;
        RECT 516.650 497.460 516.970 497.520 ;
        RECT 516.650 473.520 516.970 473.580 ;
        RECT 1331.770 473.520 1332.090 473.580 ;
        RECT 516.650 473.380 1332.090 473.520 ;
        RECT 516.650 473.320 516.970 473.380 ;
        RECT 1331.770 473.320 1332.090 473.380 ;
      LAYER via ;
        RECT 514.150 499.500 514.410 499.760 ;
        RECT 516.680 497.460 516.940 497.720 ;
        RECT 516.680 473.320 516.940 473.580 ;
        RECT 1331.800 473.320 1332.060 473.580 ;
      LAYER met2 ;
        RECT 514.170 500.000 514.450 504.000 ;
        RECT 514.210 499.790 514.350 500.000 ;
        RECT 514.150 499.470 514.410 499.790 ;
        RECT 516.680 497.430 516.940 497.750 ;
        RECT 516.740 473.610 516.880 497.430 ;
        RECT 516.680 473.290 516.940 473.610 ;
        RECT 1331.800 473.290 1332.060 473.610 ;
        RECT 1331.860 82.870 1332.000 473.290 ;
        RECT 1331.860 82.730 1335.680 82.870 ;
        RECT 1335.540 2.400 1335.680 82.730 ;
        RECT 1335.330 -4.800 1335.890 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1345.570 16.900 1345.890 16.960 ;
        RECT 1352.010 16.900 1352.330 16.960 ;
        RECT 1345.570 16.760 1352.330 16.900 ;
        RECT 1345.570 16.700 1345.890 16.760 ;
        RECT 1352.010 16.700 1352.330 16.760 ;
      LAYER via ;
        RECT 1345.600 16.700 1345.860 16.960 ;
        RECT 1352.040 16.700 1352.300 16.960 ;
      LAYER met2 ;
        RECT 515.550 500.000 515.830 504.000 ;
        RECT 515.590 499.815 515.730 500.000 ;
        RECT 515.520 499.445 515.800 499.815 ;
        RECT 515.290 491.115 515.570 491.485 ;
        RECT 515.360 477.885 515.500 491.115 ;
        RECT 515.290 477.515 515.570 477.885 ;
        RECT 1345.590 134.795 1345.870 135.165 ;
        RECT 1345.660 16.990 1345.800 134.795 ;
        RECT 1345.600 16.670 1345.860 16.990 ;
        RECT 1352.040 16.670 1352.300 16.990 ;
        RECT 1352.100 2.400 1352.240 16.670 ;
        RECT 1351.890 -4.800 1352.450 2.400 ;
      LAYER via2 ;
        RECT 515.520 499.490 515.800 499.770 ;
        RECT 515.290 491.160 515.570 491.440 ;
        RECT 515.290 477.560 515.570 477.840 ;
        RECT 1345.590 134.840 1345.870 135.120 ;
      LAYER met3 ;
        RECT 514.550 499.610 514.930 499.620 ;
        RECT 515.495 499.610 515.825 499.795 ;
        RECT 514.550 499.465 515.825 499.610 ;
        RECT 514.550 499.310 515.810 499.465 ;
        RECT 514.550 499.300 514.930 499.310 ;
        RECT 514.550 491.450 514.930 491.460 ;
        RECT 515.265 491.450 515.595 491.465 ;
        RECT 514.550 491.150 515.595 491.450 ;
        RECT 514.550 491.140 514.930 491.150 ;
        RECT 515.265 491.135 515.595 491.150 ;
        RECT 514.550 477.850 514.930 477.860 ;
        RECT 515.265 477.850 515.595 477.865 ;
        RECT 514.550 477.550 515.595 477.850 ;
        RECT 514.550 477.540 514.930 477.550 ;
        RECT 515.265 477.535 515.595 477.550 ;
        RECT 514.550 135.130 514.930 135.140 ;
        RECT 1345.565 135.130 1345.895 135.145 ;
        RECT 514.550 134.830 1345.895 135.130 ;
        RECT 514.550 134.820 514.930 134.830 ;
        RECT 1345.565 134.815 1345.895 134.830 ;
      LAYER via3 ;
        RECT 514.580 499.300 514.900 499.620 ;
        RECT 514.580 491.140 514.900 491.460 ;
        RECT 514.580 477.540 514.900 477.860 ;
        RECT 514.580 134.820 514.900 135.140 ;
      LAYER met4 ;
        RECT 514.575 499.295 514.905 499.625 ;
        RECT 514.590 491.465 514.890 499.295 ;
        RECT 514.575 491.135 514.905 491.465 ;
        RECT 514.575 477.535 514.905 477.865 ;
        RECT 514.590 135.145 514.890 477.535 ;
        RECT 514.575 134.815 514.905 135.145 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.670 136.240 464.990 136.300 ;
        RECT 752.170 136.240 752.490 136.300 ;
        RECT 464.670 136.100 752.490 136.240 ;
        RECT 464.670 136.040 464.990 136.100 ;
        RECT 752.170 136.040 752.490 136.100 ;
      LAYER via ;
        RECT 464.700 136.040 464.960 136.300 ;
        RECT 752.200 136.040 752.460 136.300 ;
      LAYER met2 ;
        RECT 465.870 500.000 466.150 504.000 ;
        RECT 465.910 498.680 466.050 500.000 ;
        RECT 465.220 498.540 466.050 498.680 ;
        RECT 465.220 472.330 465.360 498.540 ;
        RECT 464.760 472.190 465.360 472.330 ;
        RECT 464.760 136.330 464.900 472.190 ;
        RECT 464.700 136.010 464.960 136.330 ;
        RECT 752.200 136.010 752.460 136.330 ;
        RECT 752.260 82.870 752.400 136.010 ;
        RECT 752.260 82.730 756.080 82.870 ;
        RECT 755.940 2.400 756.080 82.730 ;
        RECT 755.730 -4.800 756.290 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 516.880 498.820 517.200 499.080 ;
        RECT 516.970 498.400 517.110 498.820 ;
        RECT 516.650 498.200 517.110 498.400 ;
        RECT 516.650 498.140 516.970 498.200 ;
      LAYER via ;
        RECT 516.910 498.820 517.170 499.080 ;
        RECT 516.680 498.140 516.940 498.400 ;
      LAYER met2 ;
        RECT 516.930 500.000 517.210 504.000 ;
        RECT 516.970 499.110 517.110 500.000 ;
        RECT 516.910 498.790 517.170 499.110 ;
        RECT 516.680 498.285 516.940 498.430 ;
        RECT 516.670 497.915 516.950 498.285 ;
        RECT 1366.290 134.115 1366.570 134.485 ;
        RECT 1366.360 82.870 1366.500 134.115 ;
        RECT 1366.360 82.730 1368.800 82.870 ;
        RECT 1368.660 2.400 1368.800 82.730 ;
        RECT 1368.450 -4.800 1369.010 2.400 ;
      LAYER via2 ;
        RECT 516.670 497.960 516.950 498.240 ;
        RECT 1366.290 134.160 1366.570 134.440 ;
      LAYER met3 ;
        RECT 515.470 498.250 515.850 498.260 ;
        RECT 516.645 498.250 516.975 498.265 ;
        RECT 515.470 497.950 516.975 498.250 ;
        RECT 515.470 497.940 515.850 497.950 ;
        RECT 516.645 497.935 516.975 497.950 ;
        RECT 515.470 134.450 515.850 134.460 ;
        RECT 1366.265 134.450 1366.595 134.465 ;
        RECT 515.470 134.150 1366.595 134.450 ;
        RECT 515.470 134.140 515.850 134.150 ;
        RECT 1366.265 134.135 1366.595 134.150 ;
      LAYER via3 ;
        RECT 515.500 497.940 515.820 498.260 ;
        RECT 515.500 134.140 515.820 134.460 ;
      LAYER met4 ;
        RECT 515.495 497.935 515.825 498.265 ;
        RECT 515.510 134.465 515.810 497.935 ;
        RECT 515.495 134.135 515.825 134.465 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.260 499.160 518.580 499.420 ;
        RECT 518.350 498.000 518.490 499.160 ;
        RECT 518.120 497.860 518.490 498.000 ;
        RECT 518.120 497.720 518.260 497.860 ;
        RECT 518.030 497.460 518.350 497.720 ;
        RECT 520.330 143.380 520.650 143.440 ;
        RECT 1380.070 143.380 1380.390 143.440 ;
        RECT 520.330 143.240 1380.390 143.380 ;
        RECT 520.330 143.180 520.650 143.240 ;
        RECT 1380.070 143.180 1380.390 143.240 ;
      LAYER via ;
        RECT 518.290 499.160 518.550 499.420 ;
        RECT 518.060 497.460 518.320 497.720 ;
        RECT 520.360 143.180 520.620 143.440 ;
        RECT 1380.100 143.180 1380.360 143.440 ;
      LAYER met2 ;
        RECT 518.310 500.000 518.590 504.000 ;
        RECT 518.350 499.450 518.490 500.000 ;
        RECT 518.290 499.130 518.550 499.450 ;
        RECT 518.060 497.430 518.320 497.750 ;
        RECT 518.120 491.485 518.260 497.430 ;
        RECT 518.050 491.115 518.330 491.485 ;
        RECT 520.350 477.515 520.630 477.885 ;
        RECT 520.420 143.470 520.560 477.515 ;
        RECT 520.360 143.150 520.620 143.470 ;
        RECT 1380.100 143.150 1380.360 143.470 ;
        RECT 1380.160 82.870 1380.300 143.150 ;
        RECT 1380.160 82.730 1385.360 82.870 ;
        RECT 1385.220 2.400 1385.360 82.730 ;
        RECT 1385.010 -4.800 1385.570 2.400 ;
      LAYER via2 ;
        RECT 518.050 491.160 518.330 491.440 ;
        RECT 520.350 477.560 520.630 477.840 ;
      LAYER met3 ;
        RECT 518.025 491.460 518.355 491.465 ;
        RECT 518.025 491.450 518.610 491.460 ;
        RECT 518.025 491.150 518.810 491.450 ;
        RECT 518.025 491.140 518.610 491.150 ;
        RECT 518.025 491.135 518.355 491.140 ;
        RECT 518.230 477.850 518.610 477.860 ;
        RECT 520.325 477.850 520.655 477.865 ;
        RECT 518.230 477.550 520.655 477.850 ;
        RECT 518.230 477.540 518.610 477.550 ;
        RECT 520.325 477.535 520.655 477.550 ;
      LAYER via3 ;
        RECT 518.260 491.140 518.580 491.460 ;
        RECT 518.260 477.540 518.580 477.860 ;
      LAYER met4 ;
        RECT 518.255 491.135 518.585 491.465 ;
        RECT 518.270 477.865 518.570 491.135 ;
        RECT 518.255 477.535 518.585 477.865 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 519.640 499.500 519.960 499.760 ;
        RECT 519.730 499.360 519.870 499.500 ;
        RECT 519.730 499.220 520.100 499.360 ;
        RECT 519.960 498.400 520.100 499.220 ;
        RECT 519.870 498.140 520.190 498.400 ;
        RECT 519.870 143.040 520.190 143.100 ;
        RECT 1400.770 143.040 1401.090 143.100 ;
        RECT 519.870 142.900 1401.090 143.040 ;
        RECT 519.870 142.840 520.190 142.900 ;
        RECT 1400.770 142.840 1401.090 142.900 ;
      LAYER via ;
        RECT 519.670 499.500 519.930 499.760 ;
        RECT 519.900 498.140 520.160 498.400 ;
        RECT 519.900 142.840 520.160 143.100 ;
        RECT 1400.800 142.840 1401.060 143.100 ;
      LAYER met2 ;
        RECT 519.690 500.000 519.970 504.000 ;
        RECT 519.730 499.790 519.870 500.000 ;
        RECT 519.670 499.470 519.930 499.790 ;
        RECT 519.900 498.110 520.160 498.430 ;
        RECT 519.960 143.130 520.100 498.110 ;
        RECT 519.900 142.810 520.160 143.130 ;
        RECT 1400.800 142.810 1401.060 143.130 ;
        RECT 1400.860 17.410 1401.000 142.810 ;
        RECT 1400.860 17.270 1401.920 17.410 ;
        RECT 1401.780 2.400 1401.920 17.270 ;
        RECT 1401.570 -4.800 1402.130 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.710 432.040 522.030 432.100 ;
        RECT 1414.570 432.040 1414.890 432.100 ;
        RECT 521.710 431.900 1414.890 432.040 ;
        RECT 521.710 431.840 522.030 431.900 ;
        RECT 1414.570 431.840 1414.890 431.900 ;
      LAYER via ;
        RECT 521.740 431.840 522.000 432.100 ;
        RECT 1414.600 431.840 1414.860 432.100 ;
      LAYER met2 ;
        RECT 521.070 500.000 521.350 504.000 ;
        RECT 521.110 499.475 521.250 500.000 ;
        RECT 521.040 499.105 521.320 499.475 ;
        RECT 520.810 497.915 521.090 498.285 ;
        RECT 520.880 479.130 521.020 497.915 ;
        RECT 520.880 478.990 521.480 479.130 ;
        RECT 521.340 478.280 521.480 478.990 ;
        RECT 521.340 478.140 521.940 478.280 ;
        RECT 521.800 432.130 521.940 478.140 ;
        RECT 521.740 431.810 522.000 432.130 ;
        RECT 1414.600 431.810 1414.860 432.130 ;
        RECT 1414.660 82.870 1414.800 431.810 ;
        RECT 1414.660 82.730 1418.480 82.870 ;
        RECT 1418.340 2.400 1418.480 82.730 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 521.040 499.150 521.320 499.430 ;
        RECT 520.810 497.960 521.090 498.240 ;
      LAYER met3 ;
        RECT 521.015 499.125 521.345 499.455 ;
        RECT 521.030 498.265 521.330 499.125 ;
        RECT 520.785 497.950 521.330 498.265 ;
        RECT 520.785 497.935 521.115 497.950 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.400 499.360 522.720 499.420 ;
        RECT 522.400 499.220 523.320 499.360 ;
        RECT 522.400 499.160 522.720 499.220 ;
        RECT 523.180 499.080 523.320 499.220 ;
        RECT 523.090 498.820 523.410 499.080 ;
        RECT 1428.370 16.900 1428.690 16.960 ;
        RECT 1434.810 16.900 1435.130 16.960 ;
        RECT 1428.370 16.760 1435.130 16.900 ;
        RECT 1428.370 16.700 1428.690 16.760 ;
        RECT 1434.810 16.700 1435.130 16.760 ;
      LAYER via ;
        RECT 522.430 499.160 522.690 499.420 ;
        RECT 523.120 498.820 523.380 499.080 ;
        RECT 1428.400 16.700 1428.660 16.960 ;
        RECT 1434.840 16.700 1435.100 16.960 ;
      LAYER met2 ;
        RECT 522.450 500.000 522.730 504.000 ;
        RECT 522.490 499.450 522.630 500.000 ;
        RECT 522.430 499.130 522.690 499.450 ;
        RECT 523.120 498.790 523.380 499.110 ;
        RECT 523.180 477.885 523.320 498.790 ;
        RECT 523.110 477.515 523.390 477.885 ;
        RECT 1428.390 140.915 1428.670 141.285 ;
        RECT 1428.460 16.990 1428.600 140.915 ;
        RECT 1428.400 16.670 1428.660 16.990 ;
        RECT 1434.840 16.670 1435.100 16.990 ;
        RECT 1434.900 2.400 1435.040 16.670 ;
        RECT 1434.690 -4.800 1435.250 2.400 ;
      LAYER via2 ;
        RECT 523.110 477.560 523.390 477.840 ;
        RECT 1428.390 140.960 1428.670 141.240 ;
      LAYER met3 ;
        RECT 521.910 477.850 522.290 477.860 ;
        RECT 523.085 477.850 523.415 477.865 ;
        RECT 521.910 477.550 523.415 477.850 ;
        RECT 521.910 477.540 522.290 477.550 ;
        RECT 523.085 477.535 523.415 477.550 ;
        RECT 521.910 141.250 522.290 141.260 ;
        RECT 1428.365 141.250 1428.695 141.265 ;
        RECT 521.910 140.950 1428.695 141.250 ;
        RECT 521.910 140.940 522.290 140.950 ;
        RECT 1428.365 140.935 1428.695 140.950 ;
      LAYER via3 ;
        RECT 521.940 477.540 522.260 477.860 ;
        RECT 521.940 140.940 522.260 141.260 ;
      LAYER met4 ;
        RECT 521.935 477.535 522.265 477.865 ;
        RECT 521.950 141.265 522.250 477.535 ;
        RECT 521.935 140.935 522.265 141.265 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.010 499.360 524.330 499.420 ;
        RECT 523.640 499.220 524.330 499.360 ;
        RECT 523.640 498.740 523.780 499.220 ;
        RECT 524.010 499.160 524.330 499.220 ;
        RECT 523.550 498.480 523.870 498.740 ;
      LAYER via ;
        RECT 524.040 499.160 524.300 499.420 ;
        RECT 523.580 498.480 523.840 498.740 ;
      LAYER met2 ;
        RECT 523.830 500.000 524.110 504.000 ;
        RECT 523.870 499.530 524.010 500.000 ;
        RECT 523.870 499.450 524.240 499.530 ;
        RECT 523.870 499.390 524.300 499.450 ;
        RECT 524.040 499.130 524.300 499.390 ;
        RECT 523.580 498.450 523.840 498.770 ;
        RECT 523.640 472.445 523.780 498.450 ;
        RECT 523.570 472.075 523.850 472.445 ;
        RECT 1449.090 472.075 1449.370 472.445 ;
        RECT 1449.160 82.870 1449.300 472.075 ;
        RECT 1449.160 82.730 1451.600 82.870 ;
        RECT 1451.460 2.400 1451.600 82.730 ;
        RECT 1451.250 -4.800 1451.810 2.400 ;
      LAYER via2 ;
        RECT 523.570 472.120 523.850 472.400 ;
        RECT 1449.090 472.120 1449.370 472.400 ;
      LAYER met3 ;
        RECT 523.545 472.410 523.875 472.425 ;
        RECT 1449.065 472.410 1449.395 472.425 ;
        RECT 523.545 472.110 1449.395 472.410 ;
        RECT 523.545 472.095 523.875 472.110 ;
        RECT 1449.065 472.095 1449.395 472.110 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.160 499.360 525.480 499.420 ;
        RECT 525.020 499.160 525.480 499.360 ;
        RECT 524.010 498.340 524.330 498.400 ;
        RECT 525.020 498.340 525.160 499.160 ;
        RECT 524.010 498.200 525.160 498.340 ;
        RECT 524.010 498.140 524.330 498.200 ;
        RECT 537.350 474.540 537.670 474.600 ;
        RECT 810.590 474.540 810.910 474.600 ;
        RECT 537.350 474.400 810.910 474.540 ;
        RECT 537.350 474.340 537.670 474.400 ;
        RECT 810.590 474.340 810.910 474.400 ;
        RECT 810.590 20.640 810.910 20.700 ;
        RECT 810.590 20.500 855.670 20.640 ;
        RECT 810.590 20.440 810.910 20.500 ;
        RECT 855.530 19.960 855.670 20.500 ;
        RECT 1467.930 20.300 1468.250 20.360 ;
        RECT 1386.830 20.160 1468.250 20.300 ;
        RECT 1386.830 19.960 1386.970 20.160 ;
        RECT 1467.930 20.100 1468.250 20.160 ;
        RECT 855.530 19.820 1386.970 19.960 ;
      LAYER via ;
        RECT 525.190 499.160 525.450 499.420 ;
        RECT 524.040 498.140 524.300 498.400 ;
        RECT 537.380 474.340 537.640 474.600 ;
        RECT 810.620 474.340 810.880 474.600 ;
        RECT 810.620 20.440 810.880 20.700 ;
        RECT 1467.960 20.100 1468.220 20.360 ;
      LAYER met2 ;
        RECT 525.210 500.000 525.490 504.000 ;
        RECT 525.250 499.450 525.390 500.000 ;
        RECT 525.190 499.130 525.450 499.450 ;
        RECT 524.040 498.285 524.300 498.430 ;
        RECT 524.030 497.915 524.310 498.285 ;
        RECT 537.370 497.235 537.650 497.605 ;
        RECT 537.440 474.630 537.580 497.235 ;
        RECT 537.380 474.310 537.640 474.630 ;
        RECT 810.620 474.310 810.880 474.630 ;
        RECT 810.680 20.730 810.820 474.310 ;
        RECT 810.620 20.410 810.880 20.730 ;
        RECT 1467.960 20.070 1468.220 20.390 ;
        RECT 1468.020 2.400 1468.160 20.070 ;
        RECT 1467.810 -4.800 1468.370 2.400 ;
      LAYER via2 ;
        RECT 524.030 497.960 524.310 498.240 ;
        RECT 537.370 497.280 537.650 497.560 ;
      LAYER met3 ;
        RECT 524.005 498.250 524.335 498.265 ;
        RECT 524.005 497.950 532.370 498.250 ;
        RECT 524.005 497.935 524.335 497.950 ;
        RECT 532.070 497.570 532.370 497.950 ;
        RECT 537.345 497.570 537.675 497.585 ;
        RECT 532.070 497.270 537.675 497.570 ;
        RECT 537.345 497.255 537.675 497.270 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.540 499.500 526.860 499.760 ;
        RECT 526.630 496.980 526.770 499.500 ;
        RECT 529.990 496.980 530.310 497.040 ;
        RECT 526.630 496.840 530.310 496.980 ;
        RECT 529.990 496.780 530.310 496.840 ;
        RECT 529.990 473.180 530.310 473.240 ;
        RECT 1483.570 473.180 1483.890 473.240 ;
        RECT 529.990 473.040 1483.890 473.180 ;
        RECT 529.990 472.980 530.310 473.040 ;
        RECT 1483.570 472.980 1483.890 473.040 ;
      LAYER via ;
        RECT 526.570 499.500 526.830 499.760 ;
        RECT 530.020 496.780 530.280 497.040 ;
        RECT 530.020 472.980 530.280 473.240 ;
        RECT 1483.600 472.980 1483.860 473.240 ;
      LAYER met2 ;
        RECT 526.590 500.000 526.870 504.000 ;
        RECT 526.630 499.790 526.770 500.000 ;
        RECT 526.570 499.470 526.830 499.790 ;
        RECT 530.020 496.750 530.280 497.070 ;
        RECT 530.080 473.270 530.220 496.750 ;
        RECT 530.020 472.950 530.280 473.270 ;
        RECT 1483.600 472.950 1483.860 473.270 ;
        RECT 1483.660 17.410 1483.800 472.950 ;
        RECT 1483.660 17.270 1484.720 17.410 ;
        RECT 1484.580 2.400 1484.720 17.270 ;
        RECT 1484.370 -4.800 1484.930 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.310 141.680 526.630 141.740 ;
        RECT 1497.370 141.680 1497.690 141.740 ;
        RECT 526.310 141.540 1497.690 141.680 ;
        RECT 526.310 141.480 526.630 141.540 ;
        RECT 1497.370 141.480 1497.690 141.540 ;
      LAYER via ;
        RECT 526.340 141.480 526.600 141.740 ;
        RECT 1497.400 141.480 1497.660 141.740 ;
      LAYER met2 ;
        RECT 527.970 500.000 528.250 504.000 ;
        RECT 528.010 499.645 528.150 500.000 ;
        RECT 527.940 499.275 528.220 499.645 ;
        RECT 526.330 491.115 526.610 491.485 ;
        RECT 526.400 141.770 526.540 491.115 ;
        RECT 526.340 141.450 526.600 141.770 ;
        RECT 1497.400 141.450 1497.660 141.770 ;
        RECT 1497.460 82.870 1497.600 141.450 ;
        RECT 1497.460 82.730 1501.280 82.870 ;
        RECT 1501.140 2.400 1501.280 82.730 ;
        RECT 1500.930 -4.800 1501.490 2.400 ;
      LAYER via2 ;
        RECT 527.940 499.320 528.220 499.600 ;
        RECT 526.330 491.160 526.610 491.440 ;
      LAYER met3 ;
        RECT 526.510 499.610 526.890 499.620 ;
        RECT 527.915 499.610 528.245 499.625 ;
        RECT 526.510 499.310 528.245 499.610 ;
        RECT 526.510 499.300 526.890 499.310 ;
        RECT 527.915 499.295 528.245 499.310 ;
        RECT 526.305 491.460 526.635 491.465 ;
        RECT 526.305 491.450 526.890 491.460 ;
        RECT 526.080 491.150 526.890 491.450 ;
        RECT 526.305 491.140 526.890 491.150 ;
        RECT 526.305 491.135 526.635 491.140 ;
      LAYER via3 ;
        RECT 526.540 499.300 526.860 499.620 ;
        RECT 526.540 491.140 526.860 491.460 ;
      LAYER met4 ;
        RECT 526.535 499.295 526.865 499.625 ;
        RECT 526.550 491.465 526.850 499.295 ;
        RECT 526.535 491.135 526.865 491.465 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.150 205.260 528.470 205.320 ;
        RECT 1511.170 205.260 1511.490 205.320 ;
        RECT 528.150 205.120 1511.490 205.260 ;
        RECT 528.150 205.060 528.470 205.120 ;
        RECT 1511.170 205.060 1511.490 205.120 ;
        RECT 1511.170 16.900 1511.490 16.960 ;
        RECT 1517.610 16.900 1517.930 16.960 ;
        RECT 1511.170 16.760 1517.930 16.900 ;
        RECT 1511.170 16.700 1511.490 16.760 ;
        RECT 1517.610 16.700 1517.930 16.760 ;
      LAYER via ;
        RECT 528.180 205.060 528.440 205.320 ;
        RECT 1511.200 205.060 1511.460 205.320 ;
        RECT 1511.200 16.700 1511.460 16.960 ;
        RECT 1517.640 16.700 1517.900 16.960 ;
      LAYER met2 ;
        RECT 529.350 500.000 529.630 504.000 ;
        RECT 529.390 498.000 529.530 500.000 ;
        RECT 529.160 497.860 529.530 498.000 ;
        RECT 529.160 483.070 529.300 497.860 ;
        RECT 528.240 482.930 529.300 483.070 ;
        RECT 528.240 205.350 528.380 482.930 ;
        RECT 528.180 205.030 528.440 205.350 ;
        RECT 1511.200 205.030 1511.460 205.350 ;
        RECT 1511.260 16.990 1511.400 205.030 ;
        RECT 1511.200 16.670 1511.460 16.990 ;
        RECT 1517.640 16.670 1517.900 16.990 ;
        RECT 1517.700 2.400 1517.840 16.670 ;
        RECT 1517.490 -4.800 1518.050 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.970 16.900 766.290 16.960 ;
        RECT 772.410 16.900 772.730 16.960 ;
        RECT 765.970 16.760 772.730 16.900 ;
        RECT 765.970 16.700 766.290 16.760 ;
        RECT 772.410 16.700 772.730 16.760 ;
      LAYER via ;
        RECT 766.000 16.700 766.260 16.960 ;
        RECT 772.440 16.700 772.700 16.960 ;
      LAYER met2 ;
        RECT 467.250 500.000 467.530 504.000 ;
        RECT 467.290 498.965 467.430 500.000 ;
        RECT 467.220 498.595 467.500 498.965 ;
        RECT 765.990 473.435 766.270 473.805 ;
        RECT 766.060 16.990 766.200 473.435 ;
        RECT 766.000 16.670 766.260 16.990 ;
        RECT 772.440 16.670 772.700 16.990 ;
        RECT 772.500 2.400 772.640 16.670 ;
        RECT 772.290 -4.800 772.850 2.400 ;
      LAYER via2 ;
        RECT 467.220 498.640 467.500 498.920 ;
        RECT 765.990 473.480 766.270 473.760 ;
      LAYER met3 ;
        RECT 467.195 498.930 467.525 498.945 ;
        RECT 468.550 498.930 468.930 498.940 ;
        RECT 467.195 498.630 468.930 498.930 ;
        RECT 467.195 498.615 467.525 498.630 ;
        RECT 468.550 498.620 468.930 498.630 ;
        RECT 468.550 473.770 468.930 473.780 ;
        RECT 765.965 473.770 766.295 473.785 ;
        RECT 468.550 473.470 766.295 473.770 ;
        RECT 468.550 473.460 468.930 473.470 ;
        RECT 765.965 473.455 766.295 473.470 ;
      LAYER via3 ;
        RECT 468.580 498.620 468.900 498.940 ;
        RECT 468.580 473.460 468.900 473.780 ;
      LAYER met4 ;
        RECT 468.575 498.615 468.905 498.945 ;
        RECT 468.590 473.785 468.890 498.615 ;
        RECT 468.575 473.455 468.905 473.785 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 530.680 499.360 531.000 499.420 ;
        RECT 530.540 499.160 531.000 499.360 ;
        RECT 530.540 498.400 530.680 499.160 ;
        RECT 530.450 498.140 530.770 498.400 ;
      LAYER via ;
        RECT 530.710 499.160 530.970 499.420 ;
        RECT 530.480 498.140 530.740 498.400 ;
      LAYER met2 ;
        RECT 530.730 500.000 531.010 504.000 ;
        RECT 530.770 499.450 530.910 500.000 ;
        RECT 530.710 499.130 530.970 499.450 ;
        RECT 530.480 498.110 530.740 498.430 ;
        RECT 530.540 481.285 530.680 498.110 ;
        RECT 530.470 480.915 530.750 481.285 ;
        RECT 1531.890 147.715 1532.170 148.085 ;
        RECT 1531.960 82.870 1532.100 147.715 ;
        RECT 1531.960 82.730 1534.400 82.870 ;
        RECT 1534.260 2.400 1534.400 82.730 ;
        RECT 1534.050 -4.800 1534.610 2.400 ;
      LAYER via2 ;
        RECT 530.470 480.960 530.750 481.240 ;
        RECT 1531.890 147.760 1532.170 148.040 ;
      LAYER met3 ;
        RECT 525.590 481.250 525.970 481.260 ;
        RECT 530.445 481.250 530.775 481.265 ;
        RECT 525.590 480.950 530.775 481.250 ;
        RECT 525.590 480.940 525.970 480.950 ;
        RECT 530.445 480.935 530.775 480.950 ;
        RECT 525.590 148.050 525.970 148.060 ;
        RECT 1531.865 148.050 1532.195 148.065 ;
        RECT 525.590 147.750 1532.195 148.050 ;
        RECT 525.590 147.740 525.970 147.750 ;
        RECT 1531.865 147.735 1532.195 147.750 ;
      LAYER via3 ;
        RECT 525.620 480.940 525.940 481.260 ;
        RECT 525.620 147.740 525.940 148.060 ;
      LAYER met4 ;
        RECT 525.615 480.935 525.945 481.265 ;
        RECT 525.630 148.065 525.930 480.935 ;
        RECT 525.615 147.735 525.945 148.065 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.060 498.820 532.380 499.080 ;
        RECT 532.150 498.060 532.290 498.820 ;
        RECT 531.830 497.860 532.290 498.060 ;
        RECT 531.830 497.800 532.150 497.860 ;
        RECT 531.370 479.980 531.690 480.040 ;
        RECT 534.130 479.980 534.450 480.040 ;
        RECT 531.370 479.840 534.450 479.980 ;
        RECT 531.370 479.780 531.690 479.840 ;
        RECT 534.130 479.780 534.450 479.840 ;
        RECT 534.130 150.180 534.450 150.240 ;
        RECT 1545.670 150.180 1545.990 150.240 ;
        RECT 534.130 150.040 1545.990 150.180 ;
        RECT 534.130 149.980 534.450 150.040 ;
        RECT 1545.670 149.980 1545.990 150.040 ;
      LAYER via ;
        RECT 532.090 498.820 532.350 499.080 ;
        RECT 531.860 497.800 532.120 498.060 ;
        RECT 531.400 479.780 531.660 480.040 ;
        RECT 534.160 479.780 534.420 480.040 ;
        RECT 534.160 149.980 534.420 150.240 ;
        RECT 1545.700 149.980 1545.960 150.240 ;
      LAYER met2 ;
        RECT 532.110 500.000 532.390 504.000 ;
        RECT 532.150 499.110 532.290 500.000 ;
        RECT 532.090 498.790 532.350 499.110 ;
        RECT 531.860 497.770 532.120 498.090 ;
        RECT 531.920 481.170 532.060 497.770 ;
        RECT 531.460 481.030 532.060 481.170 ;
        RECT 531.460 480.070 531.600 481.030 ;
        RECT 531.400 479.750 531.660 480.070 ;
        RECT 534.160 479.750 534.420 480.070 ;
        RECT 534.220 150.270 534.360 479.750 ;
        RECT 534.160 149.950 534.420 150.270 ;
        RECT 1545.700 149.950 1545.960 150.270 ;
        RECT 1545.760 82.870 1545.900 149.950 ;
        RECT 1545.760 82.730 1550.960 82.870 ;
        RECT 1550.820 2.400 1550.960 82.730 ;
        RECT 1550.610 -4.800 1551.170 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 533.440 499.500 533.760 499.760 ;
        RECT 533.530 498.060 533.670 499.500 ;
        RECT 533.210 497.860 533.670 498.060 ;
        RECT 533.210 497.800 533.530 497.860 ;
        RECT 533.210 149.500 533.530 149.560 ;
        RECT 1566.830 149.500 1567.150 149.560 ;
        RECT 533.210 149.360 1567.150 149.500 ;
        RECT 533.210 149.300 533.530 149.360 ;
        RECT 1566.830 149.300 1567.150 149.360 ;
      LAYER via ;
        RECT 533.470 499.500 533.730 499.760 ;
        RECT 533.240 497.800 533.500 498.060 ;
        RECT 533.240 149.300 533.500 149.560 ;
        RECT 1566.860 149.300 1567.120 149.560 ;
      LAYER met2 ;
        RECT 533.490 500.000 533.770 504.000 ;
        RECT 533.530 499.790 533.670 500.000 ;
        RECT 533.470 499.470 533.730 499.790 ;
        RECT 533.240 497.770 533.500 498.090 ;
        RECT 533.300 149.590 533.440 497.770 ;
        RECT 533.240 149.270 533.500 149.590 ;
        RECT 1566.860 149.270 1567.120 149.590 ;
        RECT 1566.920 82.870 1567.060 149.270 ;
        RECT 1566.920 82.730 1567.520 82.870 ;
        RECT 1567.380 2.400 1567.520 82.730 ;
        RECT 1567.170 -4.800 1567.730 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.820 499.500 535.140 499.760 ;
        RECT 534.910 499.080 535.050 499.500 ;
        RECT 534.590 498.880 535.050 499.080 ;
        RECT 534.590 498.820 534.910 498.880 ;
        RECT 534.590 156.980 534.910 157.040 ;
        RECT 1580.170 156.980 1580.490 157.040 ;
        RECT 534.590 156.840 1580.490 156.980 ;
        RECT 534.590 156.780 534.910 156.840 ;
        RECT 1580.170 156.780 1580.490 156.840 ;
      LAYER via ;
        RECT 534.850 499.500 535.110 499.760 ;
        RECT 534.620 498.820 534.880 499.080 ;
        RECT 534.620 156.780 534.880 157.040 ;
        RECT 1580.200 156.780 1580.460 157.040 ;
      LAYER met2 ;
        RECT 534.870 500.000 535.150 504.000 ;
        RECT 534.910 499.790 535.050 500.000 ;
        RECT 534.850 499.470 535.110 499.790 ;
        RECT 534.620 498.790 534.880 499.110 ;
        RECT 534.680 157.070 534.820 498.790 ;
        RECT 534.620 156.750 534.880 157.070 ;
        RECT 1580.200 156.750 1580.460 157.070 ;
        RECT 1580.260 82.870 1580.400 156.750 ;
        RECT 1580.260 82.730 1584.080 82.870 ;
        RECT 1583.940 2.400 1584.080 82.730 ;
        RECT 1583.730 -4.800 1584.290 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1593.970 16.900 1594.290 16.960 ;
        RECT 1600.410 16.900 1600.730 16.960 ;
        RECT 1593.970 16.760 1600.730 16.900 ;
        RECT 1593.970 16.700 1594.290 16.760 ;
        RECT 1600.410 16.700 1600.730 16.760 ;
      LAYER via ;
        RECT 1594.000 16.700 1594.260 16.960 ;
        RECT 1600.440 16.700 1600.700 16.960 ;
      LAYER met2 ;
        RECT 536.250 500.000 536.530 504.000 ;
        RECT 536.290 498.340 536.430 500.000 ;
        RECT 536.290 498.200 536.660 498.340 ;
        RECT 536.520 481.965 536.660 498.200 ;
        RECT 536.450 481.595 536.730 481.965 ;
        RECT 1593.990 155.195 1594.270 155.565 ;
        RECT 1594.060 16.990 1594.200 155.195 ;
        RECT 1594.000 16.670 1594.260 16.990 ;
        RECT 1600.440 16.670 1600.700 16.990 ;
        RECT 1600.500 2.400 1600.640 16.670 ;
        RECT 1600.290 -4.800 1600.850 2.400 ;
      LAYER via2 ;
        RECT 536.450 481.640 536.730 481.920 ;
        RECT 1593.990 155.240 1594.270 155.520 ;
      LAYER met3 ;
        RECT 535.710 481.930 536.090 481.940 ;
        RECT 536.425 481.930 536.755 481.945 ;
        RECT 535.710 481.630 536.755 481.930 ;
        RECT 535.710 481.620 536.090 481.630 ;
        RECT 536.425 481.615 536.755 481.630 ;
        RECT 535.710 155.530 536.090 155.540 ;
        RECT 1593.965 155.530 1594.295 155.545 ;
        RECT 535.710 155.230 1594.295 155.530 ;
        RECT 535.710 155.220 536.090 155.230 ;
        RECT 1593.965 155.215 1594.295 155.230 ;
      LAYER via3 ;
        RECT 535.740 481.620 536.060 481.940 ;
        RECT 535.740 155.220 536.060 155.540 ;
      LAYER met4 ;
        RECT 535.735 481.615 536.065 481.945 ;
        RECT 535.750 155.545 536.050 481.615 ;
        RECT 535.735 155.215 536.065 155.545 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.630 500.000 537.910 504.000 ;
        RECT 537.670 499.645 537.810 500.000 ;
        RECT 537.600 499.275 537.880 499.645 ;
        RECT 537.830 498.595 538.110 498.965 ;
        RECT 537.900 481.285 538.040 498.595 ;
        RECT 537.830 480.915 538.110 481.285 ;
        RECT 1614.690 154.515 1614.970 154.885 ;
        RECT 1614.760 82.870 1614.900 154.515 ;
        RECT 1614.760 82.730 1617.200 82.870 ;
        RECT 1617.060 2.400 1617.200 82.730 ;
        RECT 1616.850 -4.800 1617.410 2.400 ;
      LAYER via2 ;
        RECT 537.600 499.320 537.880 499.600 ;
        RECT 537.830 498.640 538.110 498.920 ;
        RECT 537.830 480.960 538.110 481.240 ;
        RECT 1614.690 154.560 1614.970 154.840 ;
      LAYER met3 ;
        RECT 537.575 499.295 537.905 499.625 ;
        RECT 537.590 498.945 537.890 499.295 ;
        RECT 537.590 498.630 538.135 498.945 ;
        RECT 537.805 498.615 538.135 498.630 ;
        RECT 534.790 481.250 535.170 481.260 ;
        RECT 537.805 481.250 538.135 481.265 ;
        RECT 534.790 480.950 538.135 481.250 ;
        RECT 534.790 480.940 535.170 480.950 ;
        RECT 537.805 480.935 538.135 480.950 ;
        RECT 534.790 154.850 535.170 154.860 ;
        RECT 1614.665 154.850 1614.995 154.865 ;
        RECT 534.790 154.550 1614.995 154.850 ;
        RECT 534.790 154.540 535.170 154.550 ;
        RECT 1614.665 154.535 1614.995 154.550 ;
      LAYER via3 ;
        RECT 534.820 480.940 535.140 481.260 ;
        RECT 534.820 154.540 535.140 154.860 ;
      LAYER met4 ;
        RECT 534.815 480.935 535.145 481.265 ;
        RECT 534.830 154.865 535.130 480.935 ;
        RECT 534.815 154.535 535.145 154.865 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 470.800 539.510 470.860 ;
        RECT 542.410 470.800 542.730 470.860 ;
        RECT 539.190 470.660 542.730 470.800 ;
        RECT 539.190 470.600 539.510 470.660 ;
        RECT 542.410 470.600 542.730 470.660 ;
        RECT 541.490 450.740 541.810 450.800 ;
        RECT 542.410 450.740 542.730 450.800 ;
        RECT 541.490 450.600 542.730 450.740 ;
        RECT 541.490 450.540 541.810 450.600 ;
        RECT 542.410 450.540 542.730 450.600 ;
        RECT 541.490 156.640 541.810 156.700 ;
        RECT 1628.470 156.640 1628.790 156.700 ;
        RECT 541.490 156.500 1628.790 156.640 ;
        RECT 541.490 156.440 541.810 156.500 ;
        RECT 1628.470 156.440 1628.790 156.500 ;
      LAYER via ;
        RECT 539.220 470.600 539.480 470.860 ;
        RECT 542.440 470.600 542.700 470.860 ;
        RECT 541.520 450.540 541.780 450.800 ;
        RECT 542.440 450.540 542.700 450.800 ;
        RECT 541.520 156.440 541.780 156.700 ;
        RECT 1628.500 156.440 1628.760 156.700 ;
      LAYER met2 ;
        RECT 539.010 500.000 539.290 504.000 ;
        RECT 539.050 499.020 539.190 500.000 ;
        RECT 539.050 498.880 539.420 499.020 ;
        RECT 539.280 498.680 539.420 498.880 ;
        RECT 539.280 498.540 539.650 498.680 ;
        RECT 539.510 498.170 539.650 498.540 ;
        RECT 539.280 498.030 539.650 498.170 ;
        RECT 539.280 470.890 539.420 498.030 ;
        RECT 539.220 470.570 539.480 470.890 ;
        RECT 542.440 470.570 542.700 470.890 ;
        RECT 542.500 450.830 542.640 470.570 ;
        RECT 541.520 450.510 541.780 450.830 ;
        RECT 542.440 450.510 542.700 450.830 ;
        RECT 541.580 156.730 541.720 450.510 ;
        RECT 541.520 156.410 541.780 156.730 ;
        RECT 1628.500 156.410 1628.760 156.730 ;
        RECT 1628.560 82.870 1628.700 156.410 ;
        RECT 1628.560 82.730 1633.760 82.870 ;
        RECT 1633.620 2.400 1633.760 82.730 ;
        RECT 1633.410 -4.800 1633.970 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 540.110 467.400 540.430 467.460 ;
        RECT 1649.170 467.400 1649.490 467.460 ;
        RECT 540.110 467.260 1649.490 467.400 ;
        RECT 540.110 467.200 540.430 467.260 ;
        RECT 1649.170 467.200 1649.490 467.260 ;
      LAYER via ;
        RECT 540.140 467.200 540.400 467.460 ;
        RECT 1649.200 467.200 1649.460 467.460 ;
      LAYER met2 ;
        RECT 540.390 500.000 540.670 504.000 ;
        RECT 540.430 498.680 540.570 500.000 ;
        RECT 540.200 498.540 540.570 498.680 ;
        RECT 540.200 467.490 540.340 498.540 ;
        RECT 540.140 467.170 540.400 467.490 ;
        RECT 1649.200 467.170 1649.460 467.490 ;
        RECT 1649.260 17.410 1649.400 467.170 ;
        RECT 1649.260 17.270 1650.320 17.410 ;
        RECT 1650.180 2.400 1650.320 17.270 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.720 499.700 542.040 499.760 ;
        RECT 541.580 499.500 542.040 499.700 ;
        RECT 541.580 497.660 541.720 499.500 ;
        RECT 541.950 497.660 542.270 497.720 ;
        RECT 541.580 497.520 542.270 497.660 ;
        RECT 541.950 497.460 542.270 497.520 ;
        RECT 541.950 164.120 542.270 164.180 ;
        RECT 1662.970 164.120 1663.290 164.180 ;
        RECT 541.950 163.980 1663.290 164.120 ;
        RECT 541.950 163.920 542.270 163.980 ;
        RECT 1662.970 163.920 1663.290 163.980 ;
      LAYER via ;
        RECT 541.750 499.500 542.010 499.760 ;
        RECT 541.980 497.460 542.240 497.720 ;
        RECT 541.980 163.920 542.240 164.180 ;
        RECT 1663.000 163.920 1663.260 164.180 ;
      LAYER met2 ;
        RECT 541.770 500.000 542.050 504.000 ;
        RECT 541.810 499.790 541.950 500.000 ;
        RECT 541.750 499.470 542.010 499.790 ;
        RECT 541.980 497.430 542.240 497.750 ;
        RECT 542.040 164.210 542.180 497.430 ;
        RECT 541.980 163.890 542.240 164.210 ;
        RECT 1663.000 163.890 1663.260 164.210 ;
        RECT 1663.060 82.870 1663.200 163.890 ;
        RECT 1663.060 82.730 1666.880 82.870 ;
        RECT 1666.740 2.400 1666.880 82.730 ;
        RECT 1666.530 -4.800 1667.090 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1676.770 16.900 1677.090 16.960 ;
        RECT 1683.210 16.900 1683.530 16.960 ;
        RECT 1676.770 16.760 1683.530 16.900 ;
        RECT 1676.770 16.700 1677.090 16.760 ;
        RECT 1683.210 16.700 1683.530 16.760 ;
      LAYER via ;
        RECT 1676.800 16.700 1677.060 16.960 ;
        RECT 1683.240 16.700 1683.500 16.960 ;
      LAYER met2 ;
        RECT 543.150 500.000 543.430 504.000 ;
        RECT 543.190 499.815 543.330 500.000 ;
        RECT 543.120 499.445 543.400 499.815 ;
        RECT 1676.790 467.315 1677.070 467.685 ;
        RECT 1676.860 16.990 1677.000 467.315 ;
        RECT 1676.800 16.670 1677.060 16.990 ;
        RECT 1683.240 16.670 1683.500 16.990 ;
        RECT 1683.300 2.400 1683.440 16.670 ;
        RECT 1683.090 -4.800 1683.650 2.400 ;
      LAYER via2 ;
        RECT 543.120 499.490 543.400 499.770 ;
        RECT 1676.790 467.360 1677.070 467.640 ;
      LAYER met3 ;
        RECT 553.190 500.290 553.570 500.300 ;
        RECT 543.340 499.990 545.250 500.290 ;
        RECT 543.340 499.795 543.640 499.990 ;
        RECT 543.095 499.480 543.640 499.795 ;
        RECT 544.950 499.610 545.250 499.990 ;
        RECT 545.870 499.990 553.570 500.290 ;
        RECT 545.870 499.610 546.170 499.990 ;
        RECT 553.190 499.980 553.570 499.990 ;
        RECT 543.095 499.465 543.425 499.480 ;
        RECT 544.950 499.310 546.170 499.610 ;
        RECT 553.190 467.650 553.570 467.660 ;
        RECT 1676.765 467.650 1677.095 467.665 ;
        RECT 553.190 467.350 1677.095 467.650 ;
        RECT 553.190 467.340 553.570 467.350 ;
        RECT 1676.765 467.335 1677.095 467.350 ;
      LAYER via3 ;
        RECT 553.220 499.980 553.540 500.300 ;
        RECT 553.220 467.340 553.540 467.660 ;
      LAYER met4 ;
        RECT 553.215 499.975 553.545 500.305 ;
        RECT 553.230 467.665 553.530 499.975 ;
        RECT 553.215 467.335 553.545 467.665 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.580 500.180 468.900 500.440 ;
        RECT 466.970 498.340 467.290 498.400 ;
        RECT 468.670 498.340 468.810 500.180 ;
        RECT 466.970 498.200 468.810 498.340 ;
        RECT 466.970 498.140 467.290 498.200 ;
      LAYER via ;
        RECT 468.610 500.180 468.870 500.440 ;
        RECT 467.000 498.140 467.260 498.400 ;
      LAYER met2 ;
        RECT 468.630 500.470 468.910 504.000 ;
        RECT 468.610 500.150 468.910 500.470 ;
        RECT 468.630 500.000 468.910 500.150 ;
        RECT 467.000 498.110 467.260 498.430 ;
        RECT 467.060 491.485 467.200 498.110 ;
        RECT 466.990 491.115 467.270 491.485 ;
        RECT 786.690 210.275 786.970 210.645 ;
        RECT 786.760 82.870 786.900 210.275 ;
        RECT 786.760 82.730 789.200 82.870 ;
        RECT 789.060 2.400 789.200 82.730 ;
        RECT 788.850 -4.800 789.410 2.400 ;
      LAYER via2 ;
        RECT 466.990 491.160 467.270 491.440 ;
        RECT 786.690 210.320 786.970 210.600 ;
      LAYER met3 ;
        RECT 466.965 491.460 467.295 491.465 ;
        RECT 466.710 491.450 467.295 491.460 ;
        RECT 466.510 491.150 467.295 491.450 ;
        RECT 466.710 491.140 467.295 491.150 ;
        RECT 466.965 491.135 467.295 491.140 ;
        RECT 466.710 210.610 467.090 210.620 ;
        RECT 786.665 210.610 786.995 210.625 ;
        RECT 466.710 210.310 786.995 210.610 ;
        RECT 466.710 210.300 467.090 210.310 ;
        RECT 786.665 210.295 786.995 210.310 ;
      LAYER via3 ;
        RECT 466.740 491.140 467.060 491.460 ;
        RECT 466.740 210.300 467.060 210.620 ;
      LAYER met4 ;
        RECT 466.735 491.135 467.065 491.465 ;
        RECT 466.750 210.625 467.050 491.135 ;
        RECT 466.735 210.295 467.065 210.625 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.020 498.480 544.340 498.740 ;
        RECT 544.110 498.000 544.250 498.480 ;
        RECT 543.420 497.860 544.250 498.000 ;
        RECT 543.420 497.720 543.560 497.860 ;
        RECT 543.330 497.460 543.650 497.720 ;
      LAYER via ;
        RECT 544.050 498.480 544.310 498.740 ;
        RECT 543.360 497.460 543.620 497.720 ;
      LAYER met2 ;
        RECT 544.530 500.000 544.810 504.000 ;
        RECT 544.050 498.680 544.310 498.770 ;
        RECT 544.570 498.680 544.710 500.000 ;
        RECT 544.050 498.540 544.710 498.680 ;
        RECT 544.050 498.450 544.310 498.540 ;
        RECT 543.360 497.430 543.620 497.750 ;
        RECT 543.420 481.285 543.560 497.430 ;
        RECT 543.350 480.915 543.630 481.285 ;
        RECT 1697.490 121.195 1697.770 121.565 ;
        RECT 1697.560 82.870 1697.700 121.195 ;
        RECT 1697.560 82.730 1700.000 82.870 ;
        RECT 1699.860 2.400 1700.000 82.730 ;
        RECT 1699.650 -4.800 1700.210 2.400 ;
      LAYER via2 ;
        RECT 543.350 480.960 543.630 481.240 ;
        RECT 1697.490 121.240 1697.770 121.520 ;
      LAYER met3 ;
        RECT 543.325 481.260 543.655 481.265 ;
        RECT 543.070 481.250 543.655 481.260 ;
        RECT 542.870 480.950 543.655 481.250 ;
        RECT 543.070 480.940 543.655 480.950 ;
        RECT 543.325 480.935 543.655 480.940 ;
        RECT 543.070 121.530 543.450 121.540 ;
        RECT 1697.465 121.530 1697.795 121.545 ;
        RECT 543.070 121.230 1697.795 121.530 ;
        RECT 543.070 121.220 543.450 121.230 ;
        RECT 1697.465 121.215 1697.795 121.230 ;
      LAYER via3 ;
        RECT 543.100 480.940 543.420 481.260 ;
        RECT 543.100 121.220 543.420 121.540 ;
      LAYER met4 ;
        RECT 543.095 480.935 543.425 481.265 ;
        RECT 543.110 121.545 543.410 480.935 ;
        RECT 543.095 121.215 543.425 121.545 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.630 483.040 545.950 483.100 ;
        RECT 551.150 483.040 551.470 483.100 ;
        RECT 545.630 482.900 551.470 483.040 ;
        RECT 545.630 482.840 545.950 482.900 ;
        RECT 551.150 482.840 551.470 482.900 ;
        RECT 551.150 475.560 551.470 475.620 ;
        RECT 579.210 475.560 579.530 475.620 ;
        RECT 551.150 475.420 579.530 475.560 ;
        RECT 551.150 475.360 551.470 475.420 ;
        RECT 579.210 475.360 579.530 475.420 ;
        RECT 1711.270 472.840 1711.590 472.900 ;
        RECT 592.640 472.700 1711.590 472.840 ;
        RECT 579.210 472.500 579.530 472.560 ;
        RECT 592.640 472.500 592.780 472.700 ;
        RECT 1711.270 472.640 1711.590 472.700 ;
        RECT 579.210 472.360 592.780 472.500 ;
        RECT 579.210 472.300 579.530 472.360 ;
      LAYER via ;
        RECT 545.660 482.840 545.920 483.100 ;
        RECT 551.180 482.840 551.440 483.100 ;
        RECT 551.180 475.360 551.440 475.620 ;
        RECT 579.240 475.360 579.500 475.620 ;
        RECT 579.240 472.300 579.500 472.560 ;
        RECT 1711.300 472.640 1711.560 472.900 ;
      LAYER met2 ;
        RECT 545.910 500.000 546.190 504.000 ;
        RECT 545.950 498.850 546.090 500.000 ;
        RECT 545.720 498.710 546.090 498.850 ;
        RECT 545.720 483.130 545.860 498.710 ;
        RECT 545.660 482.810 545.920 483.130 ;
        RECT 551.180 482.810 551.440 483.130 ;
        RECT 551.240 475.650 551.380 482.810 ;
        RECT 551.180 475.330 551.440 475.650 ;
        RECT 579.240 475.330 579.500 475.650 ;
        RECT 579.300 472.590 579.440 475.330 ;
        RECT 1711.300 472.610 1711.560 472.930 ;
        RECT 579.240 472.270 579.500 472.590 ;
        RECT 1711.360 82.870 1711.500 472.610 ;
        RECT 1711.360 82.730 1716.560 82.870 ;
        RECT 1716.420 2.400 1716.560 82.730 ;
        RECT 1716.210 -4.800 1716.770 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 556.670 467.060 556.990 467.120 ;
        RECT 1731.970 467.060 1732.290 467.120 ;
        RECT 556.670 466.920 1732.290 467.060 ;
        RECT 556.670 466.860 556.990 466.920 ;
        RECT 1731.970 466.860 1732.290 466.920 ;
      LAYER via ;
        RECT 556.700 466.860 556.960 467.120 ;
        RECT 1732.000 466.860 1732.260 467.120 ;
      LAYER met2 ;
        RECT 547.290 500.000 547.570 504.000 ;
        RECT 547.330 499.645 547.470 500.000 ;
        RECT 547.260 499.275 547.540 499.645 ;
        RECT 556.690 497.235 556.970 497.605 ;
        RECT 556.760 467.150 556.900 497.235 ;
        RECT 556.700 466.830 556.960 467.150 ;
        RECT 1732.000 466.830 1732.260 467.150 ;
        RECT 1732.060 17.410 1732.200 466.830 ;
        RECT 1732.060 17.270 1733.120 17.410 ;
        RECT 1732.980 2.400 1733.120 17.270 ;
        RECT 1732.770 -4.800 1733.330 2.400 ;
      LAYER via2 ;
        RECT 547.260 499.320 547.540 499.600 ;
        RECT 556.690 497.280 556.970 497.560 ;
      LAYER met3 ;
        RECT 547.235 499.610 547.565 499.625 ;
        RECT 547.235 499.310 548.930 499.610 ;
        RECT 547.235 499.295 547.565 499.310 ;
        RECT 548.630 497.570 548.930 499.310 ;
        RECT 556.665 497.570 556.995 497.585 ;
        RECT 548.630 497.270 556.995 497.570 ;
        RECT 556.665 497.255 556.995 497.270 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 548.850 466.720 549.170 466.780 ;
        RECT 1745.770 466.720 1746.090 466.780 ;
        RECT 548.850 466.580 1746.090 466.720 ;
        RECT 548.850 466.520 549.170 466.580 ;
        RECT 1745.770 466.520 1746.090 466.580 ;
      LAYER via ;
        RECT 548.880 466.520 549.140 466.780 ;
        RECT 1745.800 466.520 1746.060 466.780 ;
      LAYER met2 ;
        RECT 548.670 500.000 548.950 504.000 ;
        RECT 548.710 498.680 548.850 500.000 ;
        RECT 548.710 498.540 549.080 498.680 ;
        RECT 548.940 466.810 549.080 498.540 ;
        RECT 548.880 466.490 549.140 466.810 ;
        RECT 1745.800 466.490 1746.060 466.810 ;
        RECT 1745.860 82.870 1746.000 466.490 ;
        RECT 1745.860 82.730 1749.680 82.870 ;
        RECT 1749.540 2.400 1749.680 82.730 ;
        RECT 1749.330 -4.800 1749.890 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 550.000 499.500 550.320 499.760 ;
        RECT 550.090 499.360 550.230 499.500 ;
        RECT 549.860 499.220 550.230 499.360 ;
        RECT 549.860 498.340 550.000 499.220 ;
        RECT 551.150 498.340 551.470 498.400 ;
        RECT 549.860 498.200 551.470 498.340 ;
        RECT 551.150 498.140 551.470 498.200 ;
        RECT 1759.570 16.900 1759.890 16.960 ;
        RECT 1766.010 16.900 1766.330 16.960 ;
        RECT 1759.570 16.760 1766.330 16.900 ;
        RECT 1759.570 16.700 1759.890 16.760 ;
        RECT 1766.010 16.700 1766.330 16.760 ;
      LAYER via ;
        RECT 550.030 499.500 550.290 499.760 ;
        RECT 551.180 498.140 551.440 498.400 ;
        RECT 1759.600 16.700 1759.860 16.960 ;
        RECT 1766.040 16.700 1766.300 16.960 ;
      LAYER met2 ;
        RECT 550.050 500.000 550.330 504.000 ;
        RECT 550.090 499.790 550.230 500.000 ;
        RECT 550.030 499.470 550.290 499.790 ;
        RECT 551.180 498.110 551.440 498.430 ;
        RECT 551.240 484.005 551.380 498.110 ;
        RECT 551.170 483.635 551.450 484.005 ;
        RECT 1759.590 120.515 1759.870 120.885 ;
        RECT 1759.660 16.990 1759.800 120.515 ;
        RECT 1759.600 16.670 1759.860 16.990 ;
        RECT 1766.040 16.670 1766.300 16.990 ;
        RECT 1766.100 2.400 1766.240 16.670 ;
        RECT 1765.890 -4.800 1766.450 2.400 ;
      LAYER via2 ;
        RECT 551.170 483.680 551.450 483.960 ;
        RECT 1759.590 120.560 1759.870 120.840 ;
      LAYER met3 ;
        RECT 546.750 483.970 547.130 483.980 ;
        RECT 551.145 483.970 551.475 483.985 ;
        RECT 546.750 483.670 551.475 483.970 ;
        RECT 546.750 483.660 547.130 483.670 ;
        RECT 551.145 483.655 551.475 483.670 ;
        RECT 546.750 120.850 547.130 120.860 ;
        RECT 1759.565 120.850 1759.895 120.865 ;
        RECT 546.750 120.550 1759.895 120.850 ;
        RECT 546.750 120.540 547.130 120.550 ;
        RECT 1759.565 120.535 1759.895 120.550 ;
      LAYER via3 ;
        RECT 546.780 483.660 547.100 483.980 ;
        RECT 546.780 120.540 547.100 120.860 ;
      LAYER met4 ;
        RECT 546.775 483.655 547.105 483.985 ;
        RECT 546.790 120.865 547.090 483.655 ;
        RECT 546.775 120.535 547.105 120.865 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 551.380 499.160 551.700 499.420 ;
        RECT 550.690 498.680 551.010 498.740 ;
        RECT 551.470 498.680 551.610 499.160 ;
        RECT 550.690 498.540 551.610 498.680 ;
        RECT 550.690 498.480 551.010 498.540 ;
      LAYER via ;
        RECT 551.410 499.160 551.670 499.420 ;
        RECT 550.720 498.480 550.980 498.740 ;
      LAYER met2 ;
        RECT 551.430 500.000 551.710 504.000 ;
        RECT 551.470 499.450 551.610 500.000 ;
        RECT 551.410 499.130 551.670 499.450 ;
        RECT 550.720 498.450 550.980 498.770 ;
        RECT 550.780 467.005 550.920 498.450 ;
        RECT 550.710 466.635 550.990 467.005 ;
        RECT 1780.290 466.635 1780.570 467.005 ;
        RECT 1780.360 82.870 1780.500 466.635 ;
        RECT 1780.360 82.730 1782.800 82.870 ;
        RECT 1782.660 2.400 1782.800 82.730 ;
        RECT 1782.450 -4.800 1783.010 2.400 ;
      LAYER via2 ;
        RECT 550.710 466.680 550.990 466.960 ;
        RECT 1780.290 466.680 1780.570 466.960 ;
      LAYER met3 ;
        RECT 550.685 466.970 551.015 466.985 ;
        RECT 1780.265 466.970 1780.595 466.985 ;
        RECT 550.685 466.670 1780.595 466.970 ;
        RECT 550.685 466.655 551.015 466.670 ;
        RECT 1780.265 466.655 1780.595 466.670 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.760 498.820 553.080 499.080 ;
        RECT 552.850 498.400 552.990 498.820 ;
        RECT 552.530 498.200 552.990 498.400 ;
        RECT 552.530 498.140 552.850 498.200 ;
        RECT 552.990 120.940 553.310 121.000 ;
        RECT 1794.070 120.940 1794.390 121.000 ;
        RECT 552.990 120.800 1794.390 120.940 ;
        RECT 552.990 120.740 553.310 120.800 ;
        RECT 1794.070 120.740 1794.390 120.800 ;
      LAYER via ;
        RECT 552.790 498.820 553.050 499.080 ;
        RECT 552.560 498.140 552.820 498.400 ;
        RECT 553.020 120.740 553.280 121.000 ;
        RECT 1794.100 120.740 1794.360 121.000 ;
      LAYER met2 ;
        RECT 552.810 500.000 553.090 504.000 ;
        RECT 552.850 499.110 552.990 500.000 ;
        RECT 552.790 498.790 553.050 499.110 ;
        RECT 552.560 498.110 552.820 498.430 ;
        RECT 552.620 485.250 552.760 498.110 ;
        RECT 552.620 485.110 553.220 485.250 ;
        RECT 553.080 121.030 553.220 485.110 ;
        RECT 553.020 120.710 553.280 121.030 ;
        RECT 1794.100 120.710 1794.360 121.030 ;
        RECT 1794.160 82.870 1794.300 120.710 ;
        RECT 1794.160 82.730 1799.360 82.870 ;
        RECT 1799.220 2.400 1799.360 82.730 ;
        RECT 1799.010 -4.800 1799.570 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.140 499.500 554.460 499.760 ;
        RECT 554.230 498.000 554.370 499.500 ;
        RECT 555.290 498.000 555.610 498.060 ;
        RECT 554.230 497.860 555.610 498.000 ;
        RECT 555.290 497.800 555.610 497.860 ;
        RECT 555.290 171.600 555.610 171.660 ;
        RECT 1815.230 171.600 1815.550 171.660 ;
        RECT 555.290 171.460 1815.550 171.600 ;
        RECT 555.290 171.400 555.610 171.460 ;
        RECT 1815.230 171.400 1815.550 171.460 ;
      LAYER via ;
        RECT 554.170 499.500 554.430 499.760 ;
        RECT 555.320 497.800 555.580 498.060 ;
        RECT 555.320 171.400 555.580 171.660 ;
        RECT 1815.260 171.400 1815.520 171.660 ;
      LAYER met2 ;
        RECT 554.190 500.000 554.470 504.000 ;
        RECT 554.230 499.790 554.370 500.000 ;
        RECT 554.170 499.470 554.430 499.790 ;
        RECT 555.320 497.770 555.580 498.090 ;
        RECT 555.380 171.690 555.520 497.770 ;
        RECT 555.320 171.370 555.580 171.690 ;
        RECT 1815.260 171.370 1815.520 171.690 ;
        RECT 1815.320 82.870 1815.460 171.370 ;
        RECT 1815.320 82.730 1815.920 82.870 ;
        RECT 1815.780 2.400 1815.920 82.730 ;
        RECT 1815.570 -4.800 1816.130 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.520 499.500 555.840 499.760 ;
        RECT 555.610 499.080 555.750 499.500 ;
        RECT 555.610 498.880 556.070 499.080 ;
        RECT 555.750 498.820 556.070 498.880 ;
        RECT 554.830 489.840 555.150 489.900 ;
        RECT 555.750 489.840 556.070 489.900 ;
        RECT 554.830 489.700 556.070 489.840 ;
        RECT 554.830 489.640 555.150 489.700 ;
        RECT 555.750 489.640 556.070 489.700 ;
        RECT 554.830 171.260 555.150 171.320 ;
        RECT 1828.570 171.260 1828.890 171.320 ;
        RECT 554.830 171.120 1828.890 171.260 ;
        RECT 554.830 171.060 555.150 171.120 ;
        RECT 1828.570 171.060 1828.890 171.120 ;
      LAYER via ;
        RECT 555.550 499.500 555.810 499.760 ;
        RECT 555.780 498.820 556.040 499.080 ;
        RECT 554.860 489.640 555.120 489.900 ;
        RECT 555.780 489.640 556.040 489.900 ;
        RECT 554.860 171.060 555.120 171.320 ;
        RECT 1828.600 171.060 1828.860 171.320 ;
      LAYER met2 ;
        RECT 555.570 500.000 555.850 504.000 ;
        RECT 555.610 499.790 555.750 500.000 ;
        RECT 555.550 499.470 555.810 499.790 ;
        RECT 555.780 498.790 556.040 499.110 ;
        RECT 555.840 489.930 555.980 498.790 ;
        RECT 554.860 489.610 555.120 489.930 ;
        RECT 555.780 489.610 556.040 489.930 ;
        RECT 554.920 171.350 555.060 489.610 ;
        RECT 554.860 171.030 555.120 171.350 ;
        RECT 1828.600 171.030 1828.860 171.350 ;
        RECT 1828.660 82.870 1828.800 171.030 ;
        RECT 1828.660 82.730 1832.480 82.870 ;
        RECT 1832.340 2.400 1832.480 82.730 ;
        RECT 1832.130 -4.800 1832.690 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1842.370 16.900 1842.690 16.960 ;
        RECT 1848.810 16.900 1849.130 16.960 ;
        RECT 1842.370 16.760 1849.130 16.900 ;
        RECT 1842.370 16.700 1842.690 16.760 ;
        RECT 1848.810 16.700 1849.130 16.760 ;
      LAYER via ;
        RECT 1842.400 16.700 1842.660 16.960 ;
        RECT 1848.840 16.700 1849.100 16.960 ;
      LAYER met2 ;
        RECT 556.950 500.000 557.230 504.000 ;
        RECT 556.990 499.815 557.130 500.000 ;
        RECT 556.920 499.445 557.200 499.815 ;
        RECT 1842.390 465.955 1842.670 466.325 ;
        RECT 1842.460 16.990 1842.600 465.955 ;
        RECT 1842.400 16.670 1842.660 16.990 ;
        RECT 1848.840 16.670 1849.100 16.990 ;
        RECT 1848.900 2.400 1849.040 16.670 ;
        RECT 1848.690 -4.800 1849.250 2.400 ;
      LAYER via2 ;
        RECT 556.920 499.490 557.200 499.770 ;
        RECT 1842.390 466.000 1842.670 466.280 ;
      LAYER met3 ;
        RECT 556.895 499.610 557.225 499.795 ;
        RECT 557.790 499.610 558.170 499.620 ;
        RECT 556.895 499.465 558.170 499.610 ;
        RECT 556.910 499.310 558.170 499.465 ;
        RECT 557.790 499.300 558.170 499.310 ;
        RECT 557.790 466.290 558.170 466.300 ;
        RECT 1842.365 466.290 1842.695 466.305 ;
        RECT 557.790 465.990 1842.695 466.290 ;
        RECT 557.790 465.980 558.170 465.990 ;
        RECT 1842.365 465.975 1842.695 465.990 ;
      LAYER via3 ;
        RECT 557.820 499.300 558.140 499.620 ;
        RECT 557.820 465.980 558.140 466.300 ;
      LAYER met4 ;
        RECT 557.815 499.295 558.145 499.625 ;
        RECT 557.830 466.305 558.130 499.295 ;
        RECT 557.815 465.975 558.145 466.305 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.960 499.500 470.280 499.760 ;
        RECT 470.050 498.060 470.190 499.500 ;
        RECT 469.730 497.860 470.190 498.060 ;
        RECT 469.730 497.800 470.050 497.860 ;
        RECT 469.730 150.860 470.050 150.920 ;
        RECT 800.470 150.860 800.790 150.920 ;
        RECT 469.730 150.720 800.790 150.860 ;
        RECT 469.730 150.660 470.050 150.720 ;
        RECT 800.470 150.660 800.790 150.720 ;
      LAYER via ;
        RECT 469.990 499.500 470.250 499.760 ;
        RECT 469.760 497.800 470.020 498.060 ;
        RECT 469.760 150.660 470.020 150.920 ;
        RECT 800.500 150.660 800.760 150.920 ;
      LAYER met2 ;
        RECT 470.010 500.000 470.290 504.000 ;
        RECT 470.050 499.790 470.190 500.000 ;
        RECT 469.990 499.470 470.250 499.790 ;
        RECT 469.760 497.770 470.020 498.090 ;
        RECT 469.820 150.950 469.960 497.770 ;
        RECT 469.760 150.630 470.020 150.950 ;
        RECT 800.500 150.630 800.760 150.950 ;
        RECT 800.560 82.870 800.700 150.630 ;
        RECT 800.560 82.730 805.760 82.870 ;
        RECT 805.620 2.400 805.760 82.730 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.280 499.160 558.600 499.420 ;
        RECT 558.370 498.400 558.510 499.160 ;
        RECT 558.050 498.200 558.510 498.400 ;
        RECT 558.050 498.140 558.370 498.200 ;
      LAYER via ;
        RECT 558.310 499.160 558.570 499.420 ;
        RECT 558.080 498.140 558.340 498.400 ;
      LAYER met2 ;
        RECT 558.330 500.000 558.610 504.000 ;
        RECT 558.370 499.450 558.510 500.000 ;
        RECT 558.310 499.130 558.570 499.450 ;
        RECT 558.080 498.110 558.340 498.430 ;
        RECT 558.140 496.925 558.280 498.110 ;
        RECT 558.070 496.555 558.350 496.925 ;
        RECT 1863.090 184.435 1863.370 184.805 ;
        RECT 1863.160 82.870 1863.300 184.435 ;
        RECT 1863.160 82.730 1865.600 82.870 ;
        RECT 1865.460 2.400 1865.600 82.730 ;
        RECT 1865.250 -4.800 1865.810 2.400 ;
      LAYER via2 ;
        RECT 558.070 496.600 558.350 496.880 ;
        RECT 1863.090 184.480 1863.370 184.760 ;
      LAYER met3 ;
        RECT 555.950 496.890 556.330 496.900 ;
        RECT 558.045 496.890 558.375 496.905 ;
        RECT 555.950 496.590 558.375 496.890 ;
        RECT 555.950 496.580 556.330 496.590 ;
        RECT 558.045 496.575 558.375 496.590 ;
        RECT 555.950 184.770 556.330 184.780 ;
        RECT 1863.065 184.770 1863.395 184.785 ;
        RECT 555.950 184.470 1863.395 184.770 ;
        RECT 555.950 184.460 556.330 184.470 ;
        RECT 1863.065 184.455 1863.395 184.470 ;
      LAYER via3 ;
        RECT 555.980 496.580 556.300 496.900 ;
        RECT 555.980 184.460 556.300 184.780 ;
      LAYER met4 ;
        RECT 555.975 496.575 556.305 496.905 ;
        RECT 555.990 184.785 556.290 496.575 ;
        RECT 555.975 184.455 556.305 184.785 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 128.760 559.750 128.820 ;
        RECT 1876.870 128.760 1877.190 128.820 ;
        RECT 559.430 128.620 1877.190 128.760 ;
        RECT 559.430 128.560 559.750 128.620 ;
        RECT 1876.870 128.560 1877.190 128.620 ;
      LAYER via ;
        RECT 559.460 128.560 559.720 128.820 ;
        RECT 1876.900 128.560 1877.160 128.820 ;
      LAYER met2 ;
        RECT 559.710 500.000 559.990 504.000 ;
        RECT 559.750 498.850 559.890 500.000 ;
        RECT 559.520 498.710 559.890 498.850 ;
        RECT 559.520 128.850 559.660 498.710 ;
        RECT 559.460 128.530 559.720 128.850 ;
        RECT 1876.900 128.530 1877.160 128.850 ;
        RECT 1876.960 82.870 1877.100 128.530 ;
        RECT 1876.960 82.730 1882.160 82.870 ;
        RECT 1882.020 2.400 1882.160 82.730 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.890 128.420 560.210 128.480 ;
        RECT 1898.030 128.420 1898.350 128.480 ;
        RECT 559.890 128.280 1898.350 128.420 ;
        RECT 559.890 128.220 560.210 128.280 ;
        RECT 1898.030 128.220 1898.350 128.280 ;
      LAYER via ;
        RECT 559.920 128.220 560.180 128.480 ;
        RECT 1898.060 128.220 1898.320 128.480 ;
      LAYER met2 ;
        RECT 561.090 500.000 561.370 504.000 ;
        RECT 561.130 498.340 561.270 500.000 ;
        RECT 560.900 498.200 561.270 498.340 ;
        RECT 560.900 472.330 561.040 498.200 ;
        RECT 559.980 472.190 561.040 472.330 ;
        RECT 559.980 128.510 560.120 472.190 ;
        RECT 559.920 128.190 560.180 128.510 ;
        RECT 1898.060 128.190 1898.320 128.510 ;
        RECT 1898.120 82.870 1898.260 128.190 ;
        RECT 1898.120 82.730 1898.720 82.870 ;
        RECT 1898.580 2.400 1898.720 82.730 ;
        RECT 1898.370 -4.800 1898.930 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.350 471.480 560.670 471.540 ;
        RECT 562.190 471.480 562.510 471.540 ;
        RECT 560.350 471.340 562.510 471.480 ;
        RECT 560.350 471.280 560.670 471.340 ;
        RECT 562.190 471.280 562.510 471.340 ;
        RECT 560.350 128.080 560.670 128.140 ;
        RECT 1911.370 128.080 1911.690 128.140 ;
        RECT 560.350 127.940 1911.690 128.080 ;
        RECT 560.350 127.880 560.670 127.940 ;
        RECT 1911.370 127.880 1911.690 127.940 ;
      LAYER via ;
        RECT 560.380 471.280 560.640 471.540 ;
        RECT 562.220 471.280 562.480 471.540 ;
        RECT 560.380 127.880 560.640 128.140 ;
        RECT 1911.400 127.880 1911.660 128.140 ;
      LAYER met2 ;
        RECT 562.470 500.000 562.750 504.000 ;
        RECT 562.510 498.340 562.650 500.000 ;
        RECT 562.280 498.200 562.650 498.340 ;
        RECT 562.280 471.570 562.420 498.200 ;
        RECT 560.380 471.250 560.640 471.570 ;
        RECT 562.220 471.250 562.480 471.570 ;
        RECT 560.440 128.170 560.580 471.250 ;
        RECT 560.380 127.850 560.640 128.170 ;
        RECT 1911.400 127.850 1911.660 128.170 ;
        RECT 1911.460 82.870 1911.600 127.850 ;
        RECT 1911.460 82.730 1915.280 82.870 ;
        RECT 1915.140 2.400 1915.280 82.730 ;
        RECT 1914.930 -4.800 1915.490 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1925.170 16.900 1925.490 16.960 ;
        RECT 1931.610 16.900 1931.930 16.960 ;
        RECT 1925.170 16.760 1931.930 16.900 ;
        RECT 1925.170 16.700 1925.490 16.760 ;
        RECT 1931.610 16.700 1931.930 16.760 ;
      LAYER via ;
        RECT 1925.200 16.700 1925.460 16.960 ;
        RECT 1931.640 16.700 1931.900 16.960 ;
      LAYER met2 ;
        RECT 563.850 500.000 564.130 504.000 ;
        RECT 563.890 499.020 564.030 500.000 ;
        RECT 563.660 498.880 564.030 499.020 ;
        RECT 563.660 484.005 563.800 498.880 ;
        RECT 563.590 483.635 563.870 484.005 ;
        RECT 1925.190 183.755 1925.470 184.125 ;
        RECT 1925.260 16.990 1925.400 183.755 ;
        RECT 1925.200 16.670 1925.460 16.990 ;
        RECT 1931.640 16.670 1931.900 16.990 ;
        RECT 1931.700 2.400 1931.840 16.670 ;
        RECT 1931.490 -4.800 1932.050 2.400 ;
      LAYER via2 ;
        RECT 563.590 483.680 563.870 483.960 ;
        RECT 1925.190 183.800 1925.470 184.080 ;
      LAYER met3 ;
        RECT 563.565 483.980 563.895 483.985 ;
        RECT 563.310 483.970 563.895 483.980 ;
        RECT 563.110 483.670 563.895 483.970 ;
        RECT 563.310 483.660 563.895 483.670 ;
        RECT 563.565 483.655 563.895 483.660 ;
        RECT 563.310 184.090 563.690 184.100 ;
        RECT 1925.165 184.090 1925.495 184.105 ;
        RECT 563.310 183.790 1925.495 184.090 ;
        RECT 563.310 183.780 563.690 183.790 ;
        RECT 1925.165 183.775 1925.495 183.790 ;
      LAYER via3 ;
        RECT 563.340 483.660 563.660 483.980 ;
        RECT 563.340 183.780 563.660 184.100 ;
      LAYER met4 ;
        RECT 563.335 483.655 563.665 483.985 ;
        RECT 563.350 184.105 563.650 483.655 ;
        RECT 563.335 183.775 563.665 184.105 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.230 500.000 565.510 504.000 ;
        RECT 565.270 498.850 565.410 500.000 ;
        RECT 565.270 498.710 565.640 498.850 ;
        RECT 565.500 496.870 565.640 498.710 ;
        RECT 565.040 496.730 565.640 496.870 ;
        RECT 565.040 485.365 565.180 496.730 ;
        RECT 564.970 484.995 565.250 485.365 ;
        RECT 1945.890 465.275 1946.170 465.645 ;
        RECT 1945.960 82.870 1946.100 465.275 ;
        RECT 1945.960 82.730 1948.400 82.870 ;
        RECT 1948.260 2.400 1948.400 82.730 ;
        RECT 1948.050 -4.800 1948.610 2.400 ;
      LAYER via2 ;
        RECT 564.970 485.040 565.250 485.320 ;
        RECT 1945.890 465.320 1946.170 465.600 ;
      LAYER met3 ;
        RECT 562.390 485.330 562.770 485.340 ;
        RECT 564.945 485.330 565.275 485.345 ;
        RECT 562.390 485.030 565.275 485.330 ;
        RECT 562.390 485.020 562.770 485.030 ;
        RECT 564.945 485.015 565.275 485.030 ;
        RECT 562.390 465.610 562.770 465.620 ;
        RECT 1945.865 465.610 1946.195 465.625 ;
        RECT 562.390 465.310 1946.195 465.610 ;
        RECT 562.390 465.300 562.770 465.310 ;
        RECT 1945.865 465.295 1946.195 465.310 ;
      LAYER via3 ;
        RECT 562.420 485.020 562.740 485.340 ;
        RECT 562.420 465.300 562.740 465.620 ;
      LAYER met4 ;
        RECT 562.415 485.015 562.745 485.345 ;
        RECT 562.430 465.625 562.730 485.015 ;
        RECT 562.415 465.295 562.745 465.625 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.850 466.040 572.170 466.100 ;
        RECT 1959.670 466.040 1959.990 466.100 ;
        RECT 571.850 465.900 1959.990 466.040 ;
        RECT 571.850 465.840 572.170 465.900 ;
        RECT 1959.670 465.840 1959.990 465.900 ;
      LAYER via ;
        RECT 571.880 465.840 572.140 466.100 ;
        RECT 1959.700 465.840 1959.960 466.100 ;
      LAYER met2 ;
        RECT 566.610 500.000 566.890 504.000 ;
        RECT 566.650 499.645 566.790 500.000 ;
        RECT 566.580 499.275 566.860 499.645 ;
        RECT 569.570 497.235 569.850 497.605 ;
        RECT 569.640 488.085 569.780 497.235 ;
        RECT 569.570 487.715 569.850 488.085 ;
        RECT 571.870 483.635 572.150 484.005 ;
        RECT 571.940 466.130 572.080 483.635 ;
        RECT 571.880 465.810 572.140 466.130 ;
        RECT 1959.700 465.810 1959.960 466.130 ;
        RECT 1959.760 82.870 1959.900 465.810 ;
        RECT 1959.760 82.730 1964.960 82.870 ;
        RECT 1964.820 2.400 1964.960 82.730 ;
        RECT 1964.610 -4.800 1965.170 2.400 ;
      LAYER via2 ;
        RECT 566.580 499.320 566.860 499.600 ;
        RECT 569.570 497.280 569.850 497.560 ;
        RECT 569.570 487.760 569.850 488.040 ;
        RECT 571.870 483.680 572.150 483.960 ;
      LAYER met3 ;
        RECT 566.555 499.610 566.885 499.625 ;
        RECT 566.555 499.310 569.170 499.610 ;
        RECT 566.555 499.295 566.885 499.310 ;
        RECT 568.870 497.570 569.170 499.310 ;
        RECT 569.545 497.570 569.875 497.585 ;
        RECT 568.870 497.270 569.875 497.570 ;
        RECT 569.545 497.255 569.875 497.270 ;
        RECT 569.545 488.050 569.875 488.065 ;
        RECT 569.545 487.750 572.850 488.050 ;
        RECT 569.545 487.735 569.875 487.750 ;
        RECT 571.845 483.970 572.175 483.985 ;
        RECT 572.550 483.970 572.850 487.750 ;
        RECT 571.845 483.670 572.850 483.970 ;
        RECT 571.845 483.655 572.175 483.670 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.250 127.740 567.570 127.800 ;
        RECT 1980.370 127.740 1980.690 127.800 ;
        RECT 567.250 127.600 1980.690 127.740 ;
        RECT 567.250 127.540 567.570 127.600 ;
        RECT 1980.370 127.540 1980.690 127.600 ;
      LAYER via ;
        RECT 567.280 127.540 567.540 127.800 ;
        RECT 1980.400 127.540 1980.660 127.800 ;
      LAYER met2 ;
        RECT 567.990 500.000 568.270 504.000 ;
        RECT 568.030 498.850 568.170 500.000 ;
        RECT 567.800 498.710 568.170 498.850 ;
        RECT 567.800 473.010 567.940 498.710 ;
        RECT 567.340 472.870 567.940 473.010 ;
        RECT 567.340 127.830 567.480 472.870 ;
        RECT 567.280 127.510 567.540 127.830 ;
        RECT 1980.400 127.510 1980.660 127.830 ;
        RECT 1980.460 17.410 1980.600 127.510 ;
        RECT 1980.460 17.270 1981.520 17.410 ;
        RECT 1981.380 2.400 1981.520 17.270 ;
        RECT 1981.170 -4.800 1981.730 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 569.320 500.040 569.640 500.100 ;
        RECT 569.320 499.900 572.540 500.040 ;
        RECT 569.320 499.840 569.640 499.900 ;
        RECT 572.400 497.380 572.540 499.900 ;
        RECT 572.310 497.120 572.630 497.380 ;
        RECT 1994.170 472.500 1994.490 472.560 ;
        RECT 593.330 472.360 1994.490 472.500 ;
        RECT 572.310 471.480 572.630 471.540 ;
        RECT 593.330 471.480 593.470 472.360 ;
        RECT 1994.170 472.300 1994.490 472.360 ;
        RECT 572.310 471.340 593.470 471.480 ;
        RECT 572.310 471.280 572.630 471.340 ;
      LAYER via ;
        RECT 569.350 499.840 569.610 500.100 ;
        RECT 572.340 497.120 572.600 497.380 ;
        RECT 572.340 471.280 572.600 471.540 ;
        RECT 1994.200 472.300 1994.460 472.560 ;
      LAYER met2 ;
        RECT 569.370 500.130 569.650 504.000 ;
        RECT 569.350 500.000 569.650 500.130 ;
        RECT 569.350 499.810 569.610 500.000 ;
        RECT 572.340 497.090 572.600 497.410 ;
        RECT 572.400 471.570 572.540 497.090 ;
        RECT 1994.200 472.270 1994.460 472.590 ;
        RECT 572.340 471.250 572.600 471.570 ;
        RECT 1994.260 82.870 1994.400 472.270 ;
        RECT 1994.260 82.730 1998.080 82.870 ;
        RECT 1997.940 2.400 1998.080 82.730 ;
        RECT 1997.730 -4.800 1998.290 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 570.700 499.500 571.020 499.760 ;
        RECT 570.790 498.680 570.930 499.500 ;
        RECT 569.180 498.540 570.930 498.680 ;
        RECT 569.180 498.400 569.320 498.540 ;
        RECT 569.090 498.140 569.410 498.400 ;
        RECT 565.410 489.840 565.730 489.900 ;
        RECT 569.090 489.840 569.410 489.900 ;
        RECT 565.410 489.700 569.410 489.840 ;
        RECT 565.410 489.640 565.730 489.700 ;
        RECT 569.090 489.640 569.410 489.700 ;
        RECT 565.410 484.060 565.730 484.120 ;
        RECT 574.610 484.060 574.930 484.120 ;
        RECT 565.410 483.920 574.930 484.060 ;
        RECT 565.410 483.860 565.730 483.920 ;
        RECT 574.610 483.860 574.930 483.920 ;
        RECT 574.610 480.660 574.930 480.720 ;
        RECT 578.750 480.660 579.070 480.720 ;
        RECT 574.610 480.520 579.070 480.660 ;
        RECT 574.610 480.460 574.930 480.520 ;
        RECT 578.750 480.460 579.070 480.520 ;
        RECT 578.750 465.700 579.070 465.760 ;
        RECT 2007.970 465.700 2008.290 465.760 ;
        RECT 578.750 465.560 2008.290 465.700 ;
        RECT 578.750 465.500 579.070 465.560 ;
        RECT 2007.970 465.500 2008.290 465.560 ;
        RECT 2007.970 16.900 2008.290 16.960 ;
        RECT 2014.410 16.900 2014.730 16.960 ;
        RECT 2007.970 16.760 2014.730 16.900 ;
        RECT 2007.970 16.700 2008.290 16.760 ;
        RECT 2014.410 16.700 2014.730 16.760 ;
      LAYER via ;
        RECT 570.730 499.500 570.990 499.760 ;
        RECT 569.120 498.140 569.380 498.400 ;
        RECT 565.440 489.640 565.700 489.900 ;
        RECT 569.120 489.640 569.380 489.900 ;
        RECT 565.440 483.860 565.700 484.120 ;
        RECT 574.640 483.860 574.900 484.120 ;
        RECT 574.640 480.460 574.900 480.720 ;
        RECT 578.780 480.460 579.040 480.720 ;
        RECT 578.780 465.500 579.040 465.760 ;
        RECT 2008.000 465.500 2008.260 465.760 ;
        RECT 2008.000 16.700 2008.260 16.960 ;
        RECT 2014.440 16.700 2014.700 16.960 ;
      LAYER met2 ;
        RECT 570.750 500.000 571.030 504.000 ;
        RECT 570.790 499.790 570.930 500.000 ;
        RECT 570.730 499.470 570.990 499.790 ;
        RECT 569.120 498.110 569.380 498.430 ;
        RECT 569.180 489.930 569.320 498.110 ;
        RECT 565.440 489.610 565.700 489.930 ;
        RECT 569.120 489.610 569.380 489.930 ;
        RECT 565.500 484.150 565.640 489.610 ;
        RECT 565.440 483.830 565.700 484.150 ;
        RECT 574.640 483.830 574.900 484.150 ;
        RECT 574.700 480.750 574.840 483.830 ;
        RECT 574.640 480.430 574.900 480.750 ;
        RECT 578.780 480.430 579.040 480.750 ;
        RECT 578.840 465.790 578.980 480.430 ;
        RECT 578.780 465.470 579.040 465.790 ;
        RECT 2008.000 465.470 2008.260 465.790 ;
        RECT 2008.060 16.990 2008.200 465.470 ;
        RECT 2008.000 16.670 2008.260 16.990 ;
        RECT 2014.440 16.670 2014.700 16.990 ;
        RECT 2014.500 2.400 2014.640 16.670 ;
        RECT 2014.290 -4.800 2014.850 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 471.570 425.920 471.890 425.980 ;
        RECT 821.170 425.920 821.490 425.980 ;
        RECT 471.570 425.780 821.490 425.920 ;
        RECT 471.570 425.720 471.890 425.780 ;
        RECT 821.170 425.720 821.490 425.780 ;
      LAYER via ;
        RECT 471.600 425.720 471.860 425.980 ;
        RECT 821.200 425.720 821.460 425.980 ;
      LAYER met2 ;
        RECT 471.390 500.000 471.670 504.000 ;
        RECT 471.430 498.680 471.570 500.000 ;
        RECT 471.430 498.540 471.800 498.680 ;
        RECT 471.660 426.010 471.800 498.540 ;
        RECT 471.600 425.690 471.860 426.010 ;
        RECT 821.200 425.690 821.460 426.010 ;
        RECT 821.260 17.410 821.400 425.690 ;
        RECT 821.260 17.270 822.320 17.410 ;
        RECT 822.180 2.400 822.320 17.270 ;
        RECT 821.970 -4.800 822.530 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.130 500.000 572.410 504.000 ;
        RECT 572.170 498.680 572.310 500.000 ;
        RECT 572.170 498.540 572.540 498.680 ;
        RECT 572.400 498.000 572.540 498.540 ;
        RECT 571.940 497.860 572.540 498.000 ;
        RECT 571.940 484.685 572.080 497.860 ;
        RECT 571.870 484.315 572.150 484.685 ;
        RECT 2028.690 168.795 2028.970 169.165 ;
        RECT 2028.760 82.870 2028.900 168.795 ;
        RECT 2028.760 82.730 2031.200 82.870 ;
        RECT 2031.060 2.400 2031.200 82.730 ;
        RECT 2030.850 -4.800 2031.410 2.400 ;
      LAYER via2 ;
        RECT 571.870 484.360 572.150 484.640 ;
        RECT 2028.690 168.840 2028.970 169.120 ;
      LAYER met3 ;
        RECT 567.910 484.650 568.290 484.660 ;
        RECT 571.845 484.650 572.175 484.665 ;
        RECT 567.910 484.350 572.175 484.650 ;
        RECT 567.910 484.340 568.290 484.350 ;
        RECT 571.845 484.335 572.175 484.350 ;
        RECT 567.910 169.130 568.290 169.140 ;
        RECT 2028.665 169.130 2028.995 169.145 ;
        RECT 567.910 168.830 2028.995 169.130 ;
        RECT 567.910 168.820 568.290 168.830 ;
        RECT 2028.665 168.815 2028.995 168.830 ;
      LAYER via3 ;
        RECT 567.940 484.340 568.260 484.660 ;
        RECT 567.940 168.820 568.260 169.140 ;
      LAYER met4 ;
        RECT 567.935 484.335 568.265 484.665 ;
        RECT 567.950 169.145 568.250 484.335 ;
        RECT 567.935 168.815 568.265 169.145 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.550 500.240 579.210 500.380 ;
        RECT 573.550 499.760 573.690 500.240 ;
        RECT 573.460 499.500 573.780 499.760 ;
        RECT 579.070 497.720 579.210 500.240 ;
        RECT 579.070 497.520 579.530 497.720 ;
        RECT 579.210 497.460 579.530 497.520 ;
        RECT 579.210 476.920 579.530 476.980 ;
        RECT 590.710 476.920 591.030 476.980 ;
        RECT 579.210 476.780 591.030 476.920 ;
        RECT 579.210 476.720 579.530 476.780 ;
        RECT 590.710 476.720 591.030 476.780 ;
        RECT 591.170 182.820 591.490 182.880 ;
        RECT 2042.470 182.820 2042.790 182.880 ;
        RECT 591.170 182.680 2042.790 182.820 ;
        RECT 591.170 182.620 591.490 182.680 ;
        RECT 2042.470 182.620 2042.790 182.680 ;
      LAYER via ;
        RECT 573.490 499.500 573.750 499.760 ;
        RECT 579.240 497.460 579.500 497.720 ;
        RECT 579.240 476.720 579.500 476.980 ;
        RECT 590.740 476.720 591.000 476.980 ;
        RECT 591.200 182.620 591.460 182.880 ;
        RECT 2042.500 182.620 2042.760 182.880 ;
      LAYER met2 ;
        RECT 573.510 500.000 573.790 504.000 ;
        RECT 573.550 499.790 573.690 500.000 ;
        RECT 573.490 499.470 573.750 499.790 ;
        RECT 579.240 497.430 579.500 497.750 ;
        RECT 579.300 477.010 579.440 497.430 ;
        RECT 579.240 476.690 579.500 477.010 ;
        RECT 590.740 476.690 591.000 477.010 ;
        RECT 590.800 448.570 590.940 476.690 ;
        RECT 590.800 448.430 591.400 448.570 ;
        RECT 591.260 182.910 591.400 448.430 ;
        RECT 591.200 182.590 591.460 182.910 ;
        RECT 2042.500 182.590 2042.760 182.910 ;
        RECT 2042.560 82.870 2042.700 182.590 ;
        RECT 2042.560 82.730 2047.760 82.870 ;
        RECT 2047.620 2.400 2047.760 82.730 ;
        RECT 2047.410 -4.800 2047.970 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.840 499.160 575.160 499.420 ;
        RECT 574.930 498.680 575.070 499.160 ;
        RECT 573.780 498.540 575.070 498.680 ;
        RECT 573.780 496.700 573.920 498.540 ;
        RECT 573.690 496.440 574.010 496.700 ;
        RECT 574.150 95.100 574.470 95.160 ;
        RECT 845.090 95.100 845.410 95.160 ;
        RECT 574.150 94.960 845.410 95.100 ;
        RECT 574.150 94.900 574.470 94.960 ;
        RECT 845.090 94.900 845.410 94.960 ;
        RECT 845.090 19.280 845.410 19.340 ;
        RECT 2064.090 19.280 2064.410 19.340 ;
        RECT 845.090 19.140 2064.410 19.280 ;
        RECT 845.090 19.080 845.410 19.140 ;
        RECT 2064.090 19.080 2064.410 19.140 ;
      LAYER via ;
        RECT 574.870 499.160 575.130 499.420 ;
        RECT 573.720 496.440 573.980 496.700 ;
        RECT 574.180 94.900 574.440 95.160 ;
        RECT 845.120 94.900 845.380 95.160 ;
        RECT 845.120 19.080 845.380 19.340 ;
        RECT 2064.120 19.080 2064.380 19.340 ;
      LAYER met2 ;
        RECT 574.890 500.000 575.170 504.000 ;
        RECT 574.930 499.450 575.070 500.000 ;
        RECT 574.870 499.130 575.130 499.450 ;
        RECT 573.720 496.410 573.980 496.730 ;
        RECT 573.780 475.220 573.920 496.410 ;
        RECT 573.780 475.080 574.380 475.220 ;
        RECT 574.240 95.190 574.380 475.080 ;
        RECT 574.180 94.870 574.440 95.190 ;
        RECT 845.120 94.870 845.380 95.190 ;
        RECT 845.180 19.370 845.320 94.870 ;
        RECT 845.120 19.050 845.380 19.370 ;
        RECT 2064.120 19.050 2064.380 19.370 ;
        RECT 2064.180 2.400 2064.320 19.050 ;
        RECT 2063.970 -4.800 2064.530 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.610 497.660 574.930 497.720 ;
        RECT 575.990 497.660 576.310 497.720 ;
        RECT 574.610 497.520 576.310 497.660 ;
        RECT 574.610 497.460 574.930 497.520 ;
        RECT 575.990 497.460 576.310 497.520 ;
        RECT 574.610 484.740 574.930 484.800 ;
        RECT 574.610 484.600 591.400 484.740 ;
        RECT 574.610 484.540 574.930 484.600 ;
        RECT 591.260 484.400 591.400 484.600 ;
        RECT 591.260 484.260 592.780 484.400 ;
        RECT 592.640 484.120 592.780 484.260 ;
        RECT 592.550 483.860 592.870 484.120 ;
        RECT 591.630 472.160 591.950 472.220 ;
        RECT 592.550 472.160 592.870 472.220 ;
        RECT 591.630 472.020 592.870 472.160 ;
        RECT 591.630 471.960 591.950 472.020 ;
        RECT 592.550 471.960 592.870 472.020 ;
        RECT 591.630 190.640 591.950 190.700 ;
        RECT 2076.970 190.640 2077.290 190.700 ;
        RECT 591.630 190.500 2077.290 190.640 ;
        RECT 591.630 190.440 591.950 190.500 ;
        RECT 2076.970 190.440 2077.290 190.500 ;
      LAYER via ;
        RECT 574.640 497.460 574.900 497.720 ;
        RECT 576.020 497.460 576.280 497.720 ;
        RECT 574.640 484.540 574.900 484.800 ;
        RECT 592.580 483.860 592.840 484.120 ;
        RECT 591.660 471.960 591.920 472.220 ;
        RECT 592.580 471.960 592.840 472.220 ;
        RECT 591.660 190.440 591.920 190.700 ;
        RECT 2077.000 190.440 2077.260 190.700 ;
      LAYER met2 ;
        RECT 576.270 500.000 576.550 504.000 ;
        RECT 576.310 498.850 576.450 500.000 ;
        RECT 576.080 498.710 576.450 498.850 ;
        RECT 576.080 497.750 576.220 498.710 ;
        RECT 574.640 497.430 574.900 497.750 ;
        RECT 576.020 497.430 576.280 497.750 ;
        RECT 574.700 484.830 574.840 497.430 ;
        RECT 574.640 484.510 574.900 484.830 ;
        RECT 592.580 483.830 592.840 484.150 ;
        RECT 592.640 472.250 592.780 483.830 ;
        RECT 591.660 471.930 591.920 472.250 ;
        RECT 592.580 471.930 592.840 472.250 ;
        RECT 591.720 190.730 591.860 471.930 ;
        RECT 591.660 190.410 591.920 190.730 ;
        RECT 2077.000 190.410 2077.260 190.730 ;
        RECT 2077.060 82.870 2077.200 190.410 ;
        RECT 2077.060 82.730 2080.880 82.870 ;
        RECT 2080.740 2.400 2080.880 82.730 ;
        RECT 2080.530 -4.800 2081.090 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 575.990 472.500 576.310 472.560 ;
        RECT 576.910 472.500 577.230 472.560 ;
        RECT 575.990 472.360 577.230 472.500 ;
        RECT 575.990 472.300 576.310 472.360 ;
        RECT 576.910 472.300 577.230 472.360 ;
        RECT 575.990 177.380 576.310 177.440 ;
        RECT 2090.770 177.380 2091.090 177.440 ;
        RECT 575.990 177.240 2091.090 177.380 ;
        RECT 575.990 177.180 576.310 177.240 ;
        RECT 2090.770 177.180 2091.090 177.240 ;
        RECT 2090.770 16.900 2091.090 16.960 ;
        RECT 2097.210 16.900 2097.530 16.960 ;
        RECT 2090.770 16.760 2097.530 16.900 ;
        RECT 2090.770 16.700 2091.090 16.760 ;
        RECT 2097.210 16.700 2097.530 16.760 ;
      LAYER via ;
        RECT 576.020 472.300 576.280 472.560 ;
        RECT 576.940 472.300 577.200 472.560 ;
        RECT 576.020 177.180 576.280 177.440 ;
        RECT 2090.800 177.180 2091.060 177.440 ;
        RECT 2090.800 16.700 2091.060 16.960 ;
        RECT 2097.240 16.700 2097.500 16.960 ;
      LAYER met2 ;
        RECT 577.650 500.000 577.930 504.000 ;
        RECT 577.690 498.850 577.830 500.000 ;
        RECT 576.770 498.710 577.830 498.850 ;
        RECT 576.770 498.340 576.910 498.710 ;
        RECT 576.540 498.200 576.910 498.340 ;
        RECT 576.540 473.690 576.680 498.200 ;
        RECT 576.540 473.550 577.140 473.690 ;
        RECT 577.000 472.590 577.140 473.550 ;
        RECT 576.020 472.270 576.280 472.590 ;
        RECT 576.940 472.270 577.200 472.590 ;
        RECT 576.080 177.470 576.220 472.270 ;
        RECT 576.020 177.150 576.280 177.470 ;
        RECT 2090.800 177.150 2091.060 177.470 ;
        RECT 2090.860 16.990 2091.000 177.150 ;
        RECT 2090.800 16.670 2091.060 16.990 ;
        RECT 2097.240 16.670 2097.500 16.990 ;
        RECT 2097.300 2.400 2097.440 16.670 ;
        RECT 2097.090 -4.800 2097.650 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 578.750 484.060 579.070 484.120 ;
        RECT 585.190 484.060 585.510 484.120 ;
        RECT 578.750 483.920 585.510 484.060 ;
        RECT 578.750 483.860 579.070 483.920 ;
        RECT 585.190 483.860 585.510 483.920 ;
        RECT 584.730 190.300 585.050 190.360 ;
        RECT 2111.470 190.300 2111.790 190.360 ;
        RECT 584.730 190.160 2111.790 190.300 ;
        RECT 584.730 190.100 585.050 190.160 ;
        RECT 2111.470 190.100 2111.790 190.160 ;
      LAYER via ;
        RECT 578.780 483.860 579.040 484.120 ;
        RECT 585.220 483.860 585.480 484.120 ;
        RECT 584.760 190.100 585.020 190.360 ;
        RECT 2111.500 190.100 2111.760 190.360 ;
      LAYER met2 ;
        RECT 579.030 500.000 579.310 504.000 ;
        RECT 579.070 498.170 579.210 500.000 ;
        RECT 578.840 498.030 579.210 498.170 ;
        RECT 578.840 484.150 578.980 498.030 ;
        RECT 578.780 483.830 579.040 484.150 ;
        RECT 585.220 483.830 585.480 484.150 ;
        RECT 585.280 448.570 585.420 483.830 ;
        RECT 584.820 448.430 585.420 448.570 ;
        RECT 584.820 190.390 584.960 448.430 ;
        RECT 584.760 190.070 585.020 190.390 ;
        RECT 2111.500 190.070 2111.760 190.390 ;
        RECT 2111.560 82.870 2111.700 190.070 ;
        RECT 2111.560 82.730 2114.000 82.870 ;
        RECT 2113.860 2.400 2114.000 82.730 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.360 499.500 580.680 499.760 ;
        RECT 580.450 498.740 580.590 499.500 ;
        RECT 580.450 498.540 580.910 498.740 ;
        RECT 580.590 498.480 580.910 498.540 ;
        RECT 581.050 189.960 581.370 190.020 ;
        RECT 2125.270 189.960 2125.590 190.020 ;
        RECT 581.050 189.820 2125.590 189.960 ;
        RECT 581.050 189.760 581.370 189.820 ;
        RECT 2125.270 189.760 2125.590 189.820 ;
      LAYER via ;
        RECT 580.390 499.500 580.650 499.760 ;
        RECT 580.620 498.480 580.880 498.740 ;
        RECT 581.080 189.760 581.340 190.020 ;
        RECT 2125.300 189.760 2125.560 190.020 ;
      LAYER met2 ;
        RECT 580.410 500.000 580.690 504.000 ;
        RECT 580.450 499.790 580.590 500.000 ;
        RECT 580.390 499.470 580.650 499.790 ;
        RECT 580.620 498.450 580.880 498.770 ;
        RECT 580.680 498.000 580.820 498.450 ;
        RECT 580.680 497.860 581.280 498.000 ;
        RECT 581.140 190.050 581.280 497.860 ;
        RECT 581.080 189.730 581.340 190.050 ;
        RECT 2125.300 189.730 2125.560 190.050 ;
        RECT 2125.360 82.870 2125.500 189.730 ;
        RECT 2125.360 82.730 2130.560 82.870 ;
        RECT 2130.420 2.400 2130.560 82.730 ;
        RECT 2130.210 -4.800 2130.770 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 592.090 439.520 592.410 439.580 ;
        RECT 2146.430 439.520 2146.750 439.580 ;
        RECT 592.090 439.380 2146.750 439.520 ;
        RECT 592.090 439.320 592.410 439.380 ;
        RECT 2146.430 439.320 2146.750 439.380 ;
      LAYER via ;
        RECT 592.120 439.320 592.380 439.580 ;
        RECT 2146.460 439.320 2146.720 439.580 ;
      LAYER met2 ;
        RECT 581.790 500.000 582.070 504.000 ;
        RECT 581.830 499.815 581.970 500.000 ;
        RECT 581.760 499.445 582.040 499.815 ;
        RECT 591.650 484.315 591.930 484.685 ;
        RECT 591.720 482.530 591.860 484.315 ;
        RECT 591.720 482.390 592.320 482.530 ;
        RECT 592.180 439.610 592.320 482.390 ;
        RECT 592.120 439.290 592.380 439.610 ;
        RECT 2146.460 439.290 2146.720 439.610 ;
        RECT 2146.520 82.870 2146.660 439.290 ;
        RECT 2146.520 82.730 2147.120 82.870 ;
        RECT 2146.980 2.400 2147.120 82.730 ;
        RECT 2146.770 -4.800 2147.330 2.400 ;
      LAYER via2 ;
        RECT 581.760 499.490 582.040 499.770 ;
        RECT 591.650 484.360 591.930 484.640 ;
      LAYER met3 ;
        RECT 581.735 499.620 582.065 499.795 ;
        RECT 581.710 499.610 582.090 499.620 ;
        RECT 581.710 499.310 582.350 499.610 ;
        RECT 581.710 499.300 582.090 499.310 ;
        RECT 581.710 484.650 582.090 484.660 ;
        RECT 591.625 484.650 591.955 484.665 ;
        RECT 581.710 484.350 591.955 484.650 ;
        RECT 581.710 484.340 582.090 484.350 ;
        RECT 591.625 484.335 591.955 484.350 ;
      LAYER via3 ;
        RECT 581.740 499.300 582.060 499.620 ;
        RECT 581.740 484.340 582.060 484.660 ;
      LAYER met4 ;
        RECT 581.735 499.295 582.065 499.625 ;
        RECT 581.750 484.665 582.050 499.295 ;
        RECT 581.735 484.335 582.065 484.665 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 583.120 499.500 583.440 499.760 ;
        RECT 583.210 499.020 583.350 499.500 ;
        RECT 583.210 498.880 584.500 499.020 ;
        RECT 584.360 498.400 584.500 498.880 ;
        RECT 584.270 498.140 584.590 498.400 ;
        RECT 581.510 472.160 581.830 472.220 ;
        RECT 583.810 472.160 584.130 472.220 ;
        RECT 581.510 472.020 584.130 472.160 ;
        RECT 581.510 471.960 581.830 472.020 ;
        RECT 583.810 471.960 584.130 472.020 ;
        RECT 581.510 189.620 581.830 189.680 ;
        RECT 2159.770 189.620 2160.090 189.680 ;
        RECT 581.510 189.480 2160.090 189.620 ;
        RECT 581.510 189.420 581.830 189.480 ;
        RECT 2159.770 189.420 2160.090 189.480 ;
      LAYER via ;
        RECT 583.150 499.500 583.410 499.760 ;
        RECT 584.300 498.140 584.560 498.400 ;
        RECT 581.540 471.960 581.800 472.220 ;
        RECT 583.840 471.960 584.100 472.220 ;
        RECT 581.540 189.420 581.800 189.680 ;
        RECT 2159.800 189.420 2160.060 189.680 ;
      LAYER met2 ;
        RECT 583.170 500.000 583.450 504.000 ;
        RECT 583.210 499.790 583.350 500.000 ;
        RECT 583.150 499.470 583.410 499.790 ;
        RECT 584.300 498.110 584.560 498.430 ;
        RECT 584.360 483.070 584.500 498.110 ;
        RECT 583.900 482.930 584.500 483.070 ;
        RECT 583.900 472.250 584.040 482.930 ;
        RECT 581.540 471.930 581.800 472.250 ;
        RECT 583.840 471.930 584.100 472.250 ;
        RECT 581.600 189.710 581.740 471.930 ;
        RECT 581.540 189.390 581.800 189.710 ;
        RECT 2159.800 189.390 2160.060 189.710 ;
        RECT 2159.860 82.870 2160.000 189.390 ;
        RECT 2159.860 82.730 2163.680 82.870 ;
        RECT 2163.540 2.400 2163.680 82.730 ;
        RECT 2163.330 -4.800 2163.890 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 584.730 478.960 585.050 479.020 ;
        RECT 612.330 478.960 612.650 479.020 ;
        RECT 584.730 478.820 612.650 478.960 ;
        RECT 584.730 478.760 585.050 478.820 ;
        RECT 612.330 478.760 612.650 478.820 ;
        RECT 612.330 403.820 612.650 403.880 ;
        RECT 2173.570 403.820 2173.890 403.880 ;
        RECT 612.330 403.680 2173.890 403.820 ;
        RECT 612.330 403.620 612.650 403.680 ;
        RECT 2173.570 403.620 2173.890 403.680 ;
        RECT 2173.570 16.900 2173.890 16.960 ;
        RECT 2180.010 16.900 2180.330 16.960 ;
        RECT 2173.570 16.760 2180.330 16.900 ;
        RECT 2173.570 16.700 2173.890 16.760 ;
        RECT 2180.010 16.700 2180.330 16.760 ;
      LAYER via ;
        RECT 584.760 478.760 585.020 479.020 ;
        RECT 612.360 478.760 612.620 479.020 ;
        RECT 612.360 403.620 612.620 403.880 ;
        RECT 2173.600 403.620 2173.860 403.880 ;
        RECT 2173.600 16.700 2173.860 16.960 ;
        RECT 2180.040 16.700 2180.300 16.960 ;
      LAYER met2 ;
        RECT 584.550 500.000 584.830 504.000 ;
        RECT 584.590 498.850 584.730 500.000 ;
        RECT 584.590 498.710 584.960 498.850 ;
        RECT 584.820 479.050 584.960 498.710 ;
        RECT 584.760 478.730 585.020 479.050 ;
        RECT 612.360 478.730 612.620 479.050 ;
        RECT 612.420 403.910 612.560 478.730 ;
        RECT 612.360 403.590 612.620 403.910 ;
        RECT 2173.600 403.590 2173.860 403.910 ;
        RECT 2173.660 16.990 2173.800 403.590 ;
        RECT 2173.600 16.670 2173.860 16.990 ;
        RECT 2180.040 16.670 2180.300 16.990 ;
        RECT 2180.100 2.400 2180.240 16.670 ;
        RECT 2179.890 -4.800 2180.450 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.720 499.160 473.040 499.420 ;
        RECT 472.810 498.680 472.950 499.160 ;
        RECT 474.330 498.680 474.650 498.740 ;
        RECT 472.810 498.540 474.650 498.680 ;
        RECT 474.330 498.480 474.650 498.540 ;
        RECT 644.990 483.040 645.310 483.100 ;
        RECT 641.630 482.900 645.310 483.040 ;
        RECT 474.330 482.360 474.650 482.420 ;
        RECT 641.630 482.360 641.770 482.900 ;
        RECT 644.990 482.840 645.310 482.900 ;
        RECT 474.330 482.220 641.770 482.360 ;
        RECT 474.330 482.160 474.650 482.220 ;
        RECT 644.990 19.280 645.310 19.340 ;
        RECT 820.710 19.280 821.030 19.340 ;
        RECT 644.990 19.140 821.030 19.280 ;
        RECT 644.990 19.080 645.310 19.140 ;
        RECT 820.710 19.080 821.030 19.140 ;
        RECT 820.710 16.900 821.030 16.960 ;
        RECT 838.650 16.900 838.970 16.960 ;
        RECT 820.710 16.760 838.970 16.900 ;
        RECT 820.710 16.700 821.030 16.760 ;
        RECT 838.650 16.700 838.970 16.760 ;
      LAYER via ;
        RECT 472.750 499.160 473.010 499.420 ;
        RECT 474.360 498.480 474.620 498.740 ;
        RECT 474.360 482.160 474.620 482.420 ;
        RECT 645.020 482.840 645.280 483.100 ;
        RECT 645.020 19.080 645.280 19.340 ;
        RECT 820.740 19.080 821.000 19.340 ;
        RECT 820.740 16.700 821.000 16.960 ;
        RECT 838.680 16.700 838.940 16.960 ;
      LAYER met2 ;
        RECT 472.770 500.000 473.050 504.000 ;
        RECT 472.810 499.450 472.950 500.000 ;
        RECT 472.750 499.130 473.010 499.450 ;
        RECT 474.360 498.450 474.620 498.770 ;
        RECT 474.420 482.450 474.560 498.450 ;
        RECT 645.020 482.810 645.280 483.130 ;
        RECT 474.360 482.130 474.620 482.450 ;
        RECT 645.080 19.370 645.220 482.810 ;
        RECT 645.020 19.050 645.280 19.370 ;
        RECT 820.740 19.050 821.000 19.370 ;
        RECT 820.800 16.990 820.940 19.050 ;
        RECT 820.740 16.670 821.000 16.990 ;
        RECT 838.680 16.670 838.940 16.990 ;
        RECT 838.740 2.400 838.880 16.670 ;
        RECT 838.530 -4.800 839.090 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.930 500.000 586.210 504.000 ;
        RECT 585.970 498.850 586.110 500.000 ;
        RECT 585.970 498.710 586.340 498.850 ;
        RECT 586.200 498.285 586.340 498.710 ;
        RECT 586.130 497.915 586.410 498.285 ;
        RECT 2194.290 189.875 2194.570 190.245 ;
        RECT 2194.360 82.870 2194.500 189.875 ;
        RECT 2194.360 82.730 2196.800 82.870 ;
        RECT 2196.660 2.400 2196.800 82.730 ;
        RECT 2196.450 -4.800 2197.010 2.400 ;
      LAYER via2 ;
        RECT 586.130 497.960 586.410 498.240 ;
        RECT 2194.290 189.920 2194.570 190.200 ;
      LAYER met3 ;
        RECT 583.550 498.250 583.930 498.260 ;
        RECT 586.105 498.250 586.435 498.265 ;
        RECT 583.550 497.950 586.435 498.250 ;
        RECT 583.550 497.940 583.930 497.950 ;
        RECT 586.105 497.935 586.435 497.950 ;
        RECT 583.550 190.210 583.930 190.220 ;
        RECT 2194.265 190.210 2194.595 190.225 ;
        RECT 583.550 189.910 2194.595 190.210 ;
        RECT 583.550 189.900 583.930 189.910 ;
        RECT 2194.265 189.895 2194.595 189.910 ;
      LAYER via3 ;
        RECT 583.580 497.940 583.900 498.260 ;
        RECT 583.580 189.900 583.900 190.220 ;
      LAYER met4 ;
        RECT 583.575 497.935 583.905 498.265 ;
        RECT 583.590 190.225 583.890 497.935 ;
        RECT 583.575 189.895 583.905 190.225 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.260 499.500 587.580 499.760 ;
        RECT 587.350 498.740 587.490 499.500 ;
        RECT 587.350 498.540 587.810 498.740 ;
        RECT 587.490 498.480 587.810 498.540 ;
        RECT 588.410 482.700 588.730 482.760 ;
        RECT 639.470 482.700 639.790 482.760 ;
        RECT 588.410 482.560 639.790 482.700 ;
        RECT 588.410 482.500 588.730 482.560 ;
        RECT 639.470 482.500 639.790 482.560 ;
        RECT 639.470 18.940 639.790 19.000 ;
        RECT 2213.130 18.940 2213.450 19.000 ;
        RECT 639.470 18.800 2213.450 18.940 ;
        RECT 639.470 18.740 639.790 18.800 ;
        RECT 2213.130 18.740 2213.450 18.800 ;
      LAYER via ;
        RECT 587.290 499.500 587.550 499.760 ;
        RECT 587.520 498.480 587.780 498.740 ;
        RECT 588.440 482.500 588.700 482.760 ;
        RECT 639.500 482.500 639.760 482.760 ;
        RECT 639.500 18.740 639.760 19.000 ;
        RECT 2213.160 18.740 2213.420 19.000 ;
      LAYER met2 ;
        RECT 587.310 500.000 587.590 504.000 ;
        RECT 587.350 499.790 587.490 500.000 ;
        RECT 587.290 499.470 587.550 499.790 ;
        RECT 587.520 498.450 587.780 498.770 ;
        RECT 587.580 498.170 587.720 498.450 ;
        RECT 587.580 498.030 588.180 498.170 ;
        RECT 588.040 492.050 588.180 498.030 ;
        RECT 588.040 491.910 588.640 492.050 ;
        RECT 588.500 482.790 588.640 491.910 ;
        RECT 588.440 482.470 588.700 482.790 ;
        RECT 639.500 482.470 639.760 482.790 ;
        RECT 639.560 19.030 639.700 482.470 ;
        RECT 639.500 18.710 639.760 19.030 ;
        RECT 2213.160 18.710 2213.420 19.030 ;
        RECT 2213.220 2.400 2213.360 18.710 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 588.410 498.480 588.730 498.740 ;
        RECT 588.500 497.320 588.640 498.480 ;
        RECT 591.630 497.320 591.950 497.380 ;
        RECT 588.500 497.180 591.950 497.320 ;
        RECT 591.630 497.120 591.950 497.180 ;
        RECT 593.010 459.580 593.330 459.640 ;
        RECT 2228.770 459.580 2229.090 459.640 ;
        RECT 593.010 459.440 2229.090 459.580 ;
        RECT 593.010 459.380 593.330 459.440 ;
        RECT 2228.770 459.380 2229.090 459.440 ;
      LAYER via ;
        RECT 588.440 498.480 588.700 498.740 ;
        RECT 591.660 497.120 591.920 497.380 ;
        RECT 593.040 459.380 593.300 459.640 ;
        RECT 2228.800 459.380 2229.060 459.640 ;
      LAYER met2 ;
        RECT 588.690 500.000 588.970 504.000 ;
        RECT 588.730 499.530 588.870 500.000 ;
        RECT 588.500 499.390 588.870 499.530 ;
        RECT 588.500 498.770 588.640 499.390 ;
        RECT 588.440 498.450 588.700 498.770 ;
        RECT 591.660 497.090 591.920 497.410 ;
        RECT 591.720 485.250 591.860 497.090 ;
        RECT 591.720 485.110 593.240 485.250 ;
        RECT 593.100 459.670 593.240 485.110 ;
        RECT 593.040 459.350 593.300 459.670 ;
        RECT 2228.800 459.350 2229.060 459.670 ;
        RECT 2228.860 17.410 2229.000 459.350 ;
        RECT 2228.860 17.270 2229.920 17.410 ;
        RECT 2229.780 2.400 2229.920 17.270 ;
        RECT 2229.570 -4.800 2230.130 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 590.020 499.160 590.340 499.420 ;
        RECT 590.110 498.060 590.250 499.160 ;
        RECT 589.790 497.860 590.250 498.060 ;
        RECT 589.790 497.800 590.110 497.860 ;
        RECT 589.790 489.840 590.110 489.900 ;
        RECT 645.910 489.840 646.230 489.900 ;
        RECT 589.790 489.700 646.230 489.840 ;
        RECT 589.790 489.640 590.110 489.700 ;
        RECT 645.910 489.640 646.230 489.700 ;
        RECT 645.910 265.780 646.230 265.840 ;
        RECT 2242.570 265.780 2242.890 265.840 ;
        RECT 645.910 265.640 2242.890 265.780 ;
        RECT 645.910 265.580 646.230 265.640 ;
        RECT 2242.570 265.580 2242.890 265.640 ;
      LAYER via ;
        RECT 590.050 499.160 590.310 499.420 ;
        RECT 589.820 497.800 590.080 498.060 ;
        RECT 589.820 489.640 590.080 489.900 ;
        RECT 645.940 489.640 646.200 489.900 ;
        RECT 645.940 265.580 646.200 265.840 ;
        RECT 2242.600 265.580 2242.860 265.840 ;
      LAYER met2 ;
        RECT 590.070 500.000 590.350 504.000 ;
        RECT 590.110 499.450 590.250 500.000 ;
        RECT 590.050 499.130 590.310 499.450 ;
        RECT 589.820 497.770 590.080 498.090 ;
        RECT 589.880 489.930 590.020 497.770 ;
        RECT 589.820 489.610 590.080 489.930 ;
        RECT 645.940 489.610 646.200 489.930 ;
        RECT 646.000 265.870 646.140 489.610 ;
        RECT 645.940 265.550 646.200 265.870 ;
        RECT 2242.600 265.550 2242.860 265.870 ;
        RECT 2242.660 82.870 2242.800 265.550 ;
        RECT 2242.660 82.730 2246.480 82.870 ;
        RECT 2246.340 2.400 2246.480 82.730 ;
        RECT 2246.130 -4.800 2246.690 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2256.370 16.900 2256.690 16.960 ;
        RECT 2262.810 16.900 2263.130 16.960 ;
        RECT 2256.370 16.760 2263.130 16.900 ;
        RECT 2256.370 16.700 2256.690 16.760 ;
        RECT 2262.810 16.700 2263.130 16.760 ;
      LAYER via ;
        RECT 2256.400 16.700 2256.660 16.960 ;
        RECT 2262.840 16.700 2263.100 16.960 ;
      LAYER met2 ;
        RECT 591.450 500.000 591.730 504.000 ;
        RECT 591.490 499.645 591.630 500.000 ;
        RECT 591.420 499.275 591.700 499.645 ;
        RECT 2256.390 189.195 2256.670 189.565 ;
        RECT 2256.460 16.990 2256.600 189.195 ;
        RECT 2256.400 16.670 2256.660 16.990 ;
        RECT 2262.840 16.670 2263.100 16.990 ;
        RECT 2262.900 2.400 2263.040 16.670 ;
        RECT 2262.690 -4.800 2263.250 2.400 ;
      LAYER via2 ;
        RECT 591.420 499.320 591.700 499.600 ;
        RECT 2256.390 189.240 2256.670 189.520 ;
      LAYER met3 ;
        RECT 589.070 499.610 589.450 499.620 ;
        RECT 591.395 499.610 591.725 499.625 ;
        RECT 589.070 499.310 591.725 499.610 ;
        RECT 589.070 499.300 589.450 499.310 ;
        RECT 591.395 499.295 591.725 499.310 ;
        RECT 589.070 189.530 589.450 189.540 ;
        RECT 2256.365 189.530 2256.695 189.545 ;
        RECT 589.070 189.230 2256.695 189.530 ;
        RECT 589.070 189.220 589.450 189.230 ;
        RECT 2256.365 189.215 2256.695 189.230 ;
      LAYER via3 ;
        RECT 589.100 499.300 589.420 499.620 ;
        RECT 589.100 189.220 589.420 189.540 ;
      LAYER met4 ;
        RECT 589.095 499.295 589.425 499.625 ;
        RECT 589.110 189.545 589.410 499.295 ;
        RECT 589.095 189.215 589.425 189.545 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.010 486.100 593.330 486.160 ;
        RECT 645.450 486.100 645.770 486.160 ;
        RECT 593.010 485.960 645.770 486.100 ;
        RECT 593.010 485.900 593.330 485.960 ;
        RECT 645.450 485.900 645.770 485.960 ;
        RECT 645.450 265.440 645.770 265.500 ;
        RECT 2277.070 265.440 2277.390 265.500 ;
        RECT 645.450 265.300 2277.390 265.440 ;
        RECT 645.450 265.240 645.770 265.300 ;
        RECT 2277.070 265.240 2277.390 265.300 ;
      LAYER via ;
        RECT 593.040 485.900 593.300 486.160 ;
        RECT 645.480 485.900 645.740 486.160 ;
        RECT 645.480 265.240 645.740 265.500 ;
        RECT 2277.100 265.240 2277.360 265.500 ;
      LAYER met2 ;
        RECT 592.830 500.000 593.110 504.000 ;
        RECT 592.870 498.680 593.010 500.000 ;
        RECT 592.870 498.540 593.240 498.680 ;
        RECT 593.100 486.190 593.240 498.540 ;
        RECT 593.040 485.870 593.300 486.190 ;
        RECT 645.480 485.870 645.740 486.190 ;
        RECT 645.540 265.530 645.680 485.870 ;
        RECT 645.480 265.210 645.740 265.530 ;
        RECT 2277.100 265.210 2277.360 265.530 ;
        RECT 2277.160 82.870 2277.300 265.210 ;
        RECT 2277.160 82.730 2279.600 82.870 ;
        RECT 2279.460 2.400 2279.600 82.730 ;
        RECT 2279.250 -4.800 2279.810 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 484.400 594.710 484.460 ;
        RECT 597.610 484.400 597.930 484.460 ;
        RECT 594.390 484.260 597.930 484.400 ;
        RECT 594.390 484.200 594.710 484.260 ;
        RECT 597.610 484.200 597.930 484.260 ;
        RECT 597.610 469.100 597.930 469.160 ;
        RECT 640.390 469.100 640.710 469.160 ;
        RECT 597.610 468.960 640.710 469.100 ;
        RECT 597.610 468.900 597.930 468.960 ;
        RECT 640.390 468.900 640.710 468.960 ;
        RECT 640.390 18.600 640.710 18.660 ;
        RECT 2283.510 18.600 2283.830 18.660 ;
        RECT 640.390 18.460 2283.830 18.600 ;
        RECT 640.390 18.400 640.710 18.460 ;
        RECT 2283.510 18.400 2283.830 18.460 ;
        RECT 2283.510 16.900 2283.830 16.960 ;
        RECT 2295.930 16.900 2296.250 16.960 ;
        RECT 2283.510 16.760 2296.250 16.900 ;
        RECT 2283.510 16.700 2283.830 16.760 ;
        RECT 2295.930 16.700 2296.250 16.760 ;
      LAYER via ;
        RECT 594.420 484.200 594.680 484.460 ;
        RECT 597.640 484.200 597.900 484.460 ;
        RECT 597.640 468.900 597.900 469.160 ;
        RECT 640.420 468.900 640.680 469.160 ;
        RECT 640.420 18.400 640.680 18.660 ;
        RECT 2283.540 18.400 2283.800 18.660 ;
        RECT 2283.540 16.700 2283.800 16.960 ;
        RECT 2295.960 16.700 2296.220 16.960 ;
      LAYER met2 ;
        RECT 594.210 500.000 594.490 504.000 ;
        RECT 594.250 498.850 594.390 500.000 ;
        RECT 594.250 498.710 594.620 498.850 ;
        RECT 594.480 484.490 594.620 498.710 ;
        RECT 594.420 484.170 594.680 484.490 ;
        RECT 597.640 484.170 597.900 484.490 ;
        RECT 597.700 469.190 597.840 484.170 ;
        RECT 597.640 468.870 597.900 469.190 ;
        RECT 640.420 468.870 640.680 469.190 ;
        RECT 640.480 18.690 640.620 468.870 ;
        RECT 640.420 18.370 640.680 18.690 ;
        RECT 2283.540 18.370 2283.800 18.690 ;
        RECT 2283.600 16.990 2283.740 18.370 ;
        RECT 2283.540 16.670 2283.800 16.990 ;
        RECT 2295.960 16.670 2296.220 16.990 ;
        RECT 2296.020 2.400 2296.160 16.670 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 595.770 485.760 596.090 485.820 ;
        RECT 646.370 485.760 646.690 485.820 ;
        RECT 595.770 485.620 646.690 485.760 ;
        RECT 595.770 485.560 596.090 485.620 ;
        RECT 646.370 485.560 646.690 485.620 ;
        RECT 646.370 272.580 646.690 272.640 ;
        RECT 2311.570 272.580 2311.890 272.640 ;
        RECT 646.370 272.440 2311.890 272.580 ;
        RECT 646.370 272.380 646.690 272.440 ;
        RECT 2311.570 272.380 2311.890 272.440 ;
      LAYER via ;
        RECT 595.800 485.560 596.060 485.820 ;
        RECT 646.400 485.560 646.660 485.820 ;
        RECT 646.400 272.380 646.660 272.640 ;
        RECT 2311.600 272.380 2311.860 272.640 ;
      LAYER met2 ;
        RECT 595.590 500.000 595.870 504.000 ;
        RECT 595.630 499.020 595.770 500.000 ;
        RECT 595.630 498.880 596.000 499.020 ;
        RECT 595.860 485.850 596.000 498.880 ;
        RECT 595.800 485.530 596.060 485.850 ;
        RECT 646.400 485.530 646.660 485.850 ;
        RECT 646.460 272.670 646.600 485.530 ;
        RECT 646.400 272.350 646.660 272.670 ;
        RECT 2311.600 272.350 2311.860 272.670 ;
        RECT 2311.660 17.410 2311.800 272.350 ;
        RECT 2311.660 17.270 2312.720 17.410 ;
        RECT 2312.580 2.400 2312.720 17.270 ;
        RECT 2312.370 -4.800 2312.930 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.230 203.560 596.550 203.620 ;
        RECT 2325.370 203.560 2325.690 203.620 ;
        RECT 596.230 203.420 2325.690 203.560 ;
        RECT 596.230 203.360 596.550 203.420 ;
        RECT 2325.370 203.360 2325.690 203.420 ;
      LAYER via ;
        RECT 596.260 203.360 596.520 203.620 ;
        RECT 2325.400 203.360 2325.660 203.620 ;
      LAYER met2 ;
        RECT 596.970 500.000 597.250 504.000 ;
        RECT 597.010 498.170 597.150 500.000 ;
        RECT 596.780 498.030 597.150 498.170 ;
        RECT 596.780 497.490 596.920 498.030 ;
        RECT 596.320 497.350 596.920 497.490 ;
        RECT 596.320 203.650 596.460 497.350 ;
        RECT 596.260 203.330 596.520 203.650 ;
        RECT 2325.400 203.330 2325.660 203.650 ;
        RECT 2325.460 82.870 2325.600 203.330 ;
        RECT 2325.460 82.730 2329.280 82.870 ;
        RECT 2329.140 2.400 2329.280 82.730 ;
        RECT 2328.930 -4.800 2329.490 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 598.300 499.700 598.620 499.760 ;
        RECT 598.300 499.500 598.760 499.700 ;
        RECT 598.620 499.080 598.760 499.500 ;
        RECT 598.530 498.820 598.850 499.080 ;
        RECT 1479.890 486.780 1480.210 486.840 ;
        RECT 614.260 486.640 1480.210 486.780 ;
        RECT 598.530 486.440 598.850 486.500 ;
        RECT 614.260 486.440 614.400 486.640 ;
        RECT 1479.890 486.580 1480.210 486.640 ;
        RECT 598.530 486.300 614.400 486.440 ;
        RECT 598.530 486.240 598.850 486.300 ;
        RECT 1479.890 19.960 1480.210 20.020 ;
        RECT 2345.610 19.960 2345.930 20.020 ;
        RECT 1479.890 19.820 2345.930 19.960 ;
        RECT 1479.890 19.760 1480.210 19.820 ;
        RECT 2345.610 19.760 2345.930 19.820 ;
      LAYER via ;
        RECT 598.330 499.500 598.590 499.760 ;
        RECT 598.560 498.820 598.820 499.080 ;
        RECT 598.560 486.240 598.820 486.500 ;
        RECT 1479.920 486.580 1480.180 486.840 ;
        RECT 1479.920 19.760 1480.180 20.020 ;
        RECT 2345.640 19.760 2345.900 20.020 ;
      LAYER met2 ;
        RECT 598.350 500.000 598.630 504.000 ;
        RECT 598.390 499.790 598.530 500.000 ;
        RECT 598.330 499.470 598.590 499.790 ;
        RECT 598.560 498.790 598.820 499.110 ;
        RECT 598.620 486.530 598.760 498.790 ;
        RECT 1479.920 486.550 1480.180 486.870 ;
        RECT 598.560 486.210 598.820 486.530 ;
        RECT 1479.980 20.050 1480.120 486.550 ;
        RECT 1479.920 19.730 1480.180 20.050 ;
        RECT 2345.640 19.730 2345.900 20.050 ;
        RECT 2345.700 2.400 2345.840 19.730 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 493.190 20.300 493.510 20.360 ;
        RECT 854.750 20.300 855.070 20.360 ;
        RECT 493.190 20.160 855.070 20.300 ;
        RECT 493.190 20.100 493.510 20.160 ;
        RECT 854.750 20.100 855.070 20.160 ;
      LAYER via ;
        RECT 493.220 20.100 493.480 20.360 ;
        RECT 854.780 20.100 855.040 20.360 ;
      LAYER met2 ;
        RECT 474.150 500.000 474.430 504.000 ;
        RECT 474.190 499.645 474.330 500.000 ;
        RECT 474.120 499.275 474.400 499.645 ;
        RECT 493.210 444.875 493.490 445.245 ;
        RECT 493.280 20.390 493.420 444.875 ;
        RECT 493.220 20.070 493.480 20.390 ;
        RECT 854.780 20.070 855.040 20.390 ;
        RECT 854.840 10.610 854.980 20.070 ;
        RECT 854.840 10.470 855.440 10.610 ;
        RECT 855.300 2.400 855.440 10.470 ;
        RECT 855.090 -4.800 855.650 2.400 ;
      LAYER via2 ;
        RECT 474.120 499.320 474.400 499.600 ;
        RECT 493.210 444.920 493.490 445.200 ;
      LAYER met3 ;
        RECT 472.230 499.610 472.610 499.620 ;
        RECT 474.095 499.610 474.425 499.625 ;
        RECT 472.230 499.310 474.425 499.610 ;
        RECT 472.230 499.300 472.610 499.310 ;
        RECT 474.095 499.295 474.425 499.310 ;
        RECT 472.230 445.210 472.610 445.220 ;
        RECT 493.185 445.210 493.515 445.225 ;
        RECT 472.230 444.910 493.515 445.210 ;
        RECT 472.230 444.900 472.610 444.910 ;
        RECT 493.185 444.895 493.515 444.910 ;
      LAYER via3 ;
        RECT 472.260 499.300 472.580 499.620 ;
        RECT 472.260 444.900 472.580 445.220 ;
      LAYER met4 ;
        RECT 472.255 499.295 472.585 499.625 ;
        RECT 472.270 445.225 472.570 499.295 ;
        RECT 472.255 444.895 472.585 445.225 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
        RECT 8.970 -39.820 12.070 3559.500 ;
        RECT 188.970 -39.820 192.070 3559.500 ;
        RECT 368.970 -39.820 372.070 3559.500 ;
        RECT 548.970 760.000 552.070 3559.500 ;
        RECT 421.040 510.640 422.640 736.880 ;
        RECT 574.640 510.640 576.240 736.880 ;
        RECT 548.970 -39.820 552.070 490.000 ;
        RECT 728.970 -39.820 732.070 3559.500 ;
        RECT 908.970 -39.820 912.070 3559.500 ;
        RECT 1088.970 -39.820 1092.070 3559.500 ;
        RECT 1268.970 -39.820 1272.070 3559.500 ;
        RECT 1448.970 -39.820 1452.070 3559.500 ;
        RECT 1628.970 -39.820 1632.070 3559.500 ;
        RECT 1808.970 -39.820 1812.070 3559.500 ;
        RECT 1988.970 -39.820 1992.070 3559.500 ;
        RECT 2168.970 -39.820 2172.070 3559.500 ;
        RECT 2348.970 -39.820 2352.070 3559.500 ;
        RECT 2528.970 -39.820 2532.070 3559.500 ;
        RECT 2708.970 -39.820 2712.070 3559.500 ;
        RECT 2888.970 -39.820 2892.070 3559.500 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
      LAYER via4 ;
        RECT -11.420 3524.560 -10.240 3525.740 ;
        RECT -9.820 3524.560 -8.640 3525.740 ;
        RECT -11.420 3522.960 -10.240 3524.140 ;
        RECT -9.820 3522.960 -8.640 3524.140 ;
        RECT -11.420 3436.090 -10.240 3437.270 ;
        RECT -9.820 3436.090 -8.640 3437.270 ;
        RECT -11.420 3434.490 -10.240 3435.670 ;
        RECT -9.820 3434.490 -8.640 3435.670 ;
        RECT -11.420 3256.090 -10.240 3257.270 ;
        RECT -9.820 3256.090 -8.640 3257.270 ;
        RECT -11.420 3254.490 -10.240 3255.670 ;
        RECT -9.820 3254.490 -8.640 3255.670 ;
        RECT -11.420 3076.090 -10.240 3077.270 ;
        RECT -9.820 3076.090 -8.640 3077.270 ;
        RECT -11.420 3074.490 -10.240 3075.670 ;
        RECT -9.820 3074.490 -8.640 3075.670 ;
        RECT -11.420 2896.090 -10.240 2897.270 ;
        RECT -9.820 2896.090 -8.640 2897.270 ;
        RECT -11.420 2894.490 -10.240 2895.670 ;
        RECT -9.820 2894.490 -8.640 2895.670 ;
        RECT -11.420 2716.090 -10.240 2717.270 ;
        RECT -9.820 2716.090 -8.640 2717.270 ;
        RECT -11.420 2714.490 -10.240 2715.670 ;
        RECT -9.820 2714.490 -8.640 2715.670 ;
        RECT -11.420 2536.090 -10.240 2537.270 ;
        RECT -9.820 2536.090 -8.640 2537.270 ;
        RECT -11.420 2534.490 -10.240 2535.670 ;
        RECT -9.820 2534.490 -8.640 2535.670 ;
        RECT -11.420 2356.090 -10.240 2357.270 ;
        RECT -9.820 2356.090 -8.640 2357.270 ;
        RECT -11.420 2354.490 -10.240 2355.670 ;
        RECT -9.820 2354.490 -8.640 2355.670 ;
        RECT -11.420 2176.090 -10.240 2177.270 ;
        RECT -9.820 2176.090 -8.640 2177.270 ;
        RECT -11.420 2174.490 -10.240 2175.670 ;
        RECT -9.820 2174.490 -8.640 2175.670 ;
        RECT -11.420 1996.090 -10.240 1997.270 ;
        RECT -9.820 1996.090 -8.640 1997.270 ;
        RECT -11.420 1994.490 -10.240 1995.670 ;
        RECT -9.820 1994.490 -8.640 1995.670 ;
        RECT -11.420 1816.090 -10.240 1817.270 ;
        RECT -9.820 1816.090 -8.640 1817.270 ;
        RECT -11.420 1814.490 -10.240 1815.670 ;
        RECT -9.820 1814.490 -8.640 1815.670 ;
        RECT -11.420 1636.090 -10.240 1637.270 ;
        RECT -9.820 1636.090 -8.640 1637.270 ;
        RECT -11.420 1634.490 -10.240 1635.670 ;
        RECT -9.820 1634.490 -8.640 1635.670 ;
        RECT -11.420 1456.090 -10.240 1457.270 ;
        RECT -9.820 1456.090 -8.640 1457.270 ;
        RECT -11.420 1454.490 -10.240 1455.670 ;
        RECT -9.820 1454.490 -8.640 1455.670 ;
        RECT -11.420 1276.090 -10.240 1277.270 ;
        RECT -9.820 1276.090 -8.640 1277.270 ;
        RECT -11.420 1274.490 -10.240 1275.670 ;
        RECT -9.820 1274.490 -8.640 1275.670 ;
        RECT -11.420 1096.090 -10.240 1097.270 ;
        RECT -9.820 1096.090 -8.640 1097.270 ;
        RECT -11.420 1094.490 -10.240 1095.670 ;
        RECT -9.820 1094.490 -8.640 1095.670 ;
        RECT -11.420 916.090 -10.240 917.270 ;
        RECT -9.820 916.090 -8.640 917.270 ;
        RECT -11.420 914.490 -10.240 915.670 ;
        RECT -9.820 914.490 -8.640 915.670 ;
        RECT -11.420 736.090 -10.240 737.270 ;
        RECT -9.820 736.090 -8.640 737.270 ;
        RECT -11.420 734.490 -10.240 735.670 ;
        RECT -9.820 734.490 -8.640 735.670 ;
        RECT -11.420 556.090 -10.240 557.270 ;
        RECT -9.820 556.090 -8.640 557.270 ;
        RECT -11.420 554.490 -10.240 555.670 ;
        RECT -9.820 554.490 -8.640 555.670 ;
        RECT -11.420 376.090 -10.240 377.270 ;
        RECT -9.820 376.090 -8.640 377.270 ;
        RECT -11.420 374.490 -10.240 375.670 ;
        RECT -9.820 374.490 -8.640 375.670 ;
        RECT -11.420 196.090 -10.240 197.270 ;
        RECT -9.820 196.090 -8.640 197.270 ;
        RECT -11.420 194.490 -10.240 195.670 ;
        RECT -9.820 194.490 -8.640 195.670 ;
        RECT -11.420 16.090 -10.240 17.270 ;
        RECT -9.820 16.090 -8.640 17.270 ;
        RECT -11.420 14.490 -10.240 15.670 ;
        RECT -9.820 14.490 -8.640 15.670 ;
        RECT -11.420 -4.460 -10.240 -3.280 ;
        RECT -9.820 -4.460 -8.640 -3.280 ;
        RECT -11.420 -6.060 -10.240 -4.880 ;
        RECT -9.820 -6.060 -8.640 -4.880 ;
        RECT 9.130 3524.560 10.310 3525.740 ;
        RECT 10.730 3524.560 11.910 3525.740 ;
        RECT 9.130 3522.960 10.310 3524.140 ;
        RECT 10.730 3522.960 11.910 3524.140 ;
        RECT 9.130 3436.090 10.310 3437.270 ;
        RECT 10.730 3436.090 11.910 3437.270 ;
        RECT 9.130 3434.490 10.310 3435.670 ;
        RECT 10.730 3434.490 11.910 3435.670 ;
        RECT 9.130 3256.090 10.310 3257.270 ;
        RECT 10.730 3256.090 11.910 3257.270 ;
        RECT 9.130 3254.490 10.310 3255.670 ;
        RECT 10.730 3254.490 11.910 3255.670 ;
        RECT 9.130 3076.090 10.310 3077.270 ;
        RECT 10.730 3076.090 11.910 3077.270 ;
        RECT 9.130 3074.490 10.310 3075.670 ;
        RECT 10.730 3074.490 11.910 3075.670 ;
        RECT 9.130 2896.090 10.310 2897.270 ;
        RECT 10.730 2896.090 11.910 2897.270 ;
        RECT 9.130 2894.490 10.310 2895.670 ;
        RECT 10.730 2894.490 11.910 2895.670 ;
        RECT 9.130 2716.090 10.310 2717.270 ;
        RECT 10.730 2716.090 11.910 2717.270 ;
        RECT 9.130 2714.490 10.310 2715.670 ;
        RECT 10.730 2714.490 11.910 2715.670 ;
        RECT 9.130 2536.090 10.310 2537.270 ;
        RECT 10.730 2536.090 11.910 2537.270 ;
        RECT 9.130 2534.490 10.310 2535.670 ;
        RECT 10.730 2534.490 11.910 2535.670 ;
        RECT 9.130 2356.090 10.310 2357.270 ;
        RECT 10.730 2356.090 11.910 2357.270 ;
        RECT 9.130 2354.490 10.310 2355.670 ;
        RECT 10.730 2354.490 11.910 2355.670 ;
        RECT 9.130 2176.090 10.310 2177.270 ;
        RECT 10.730 2176.090 11.910 2177.270 ;
        RECT 9.130 2174.490 10.310 2175.670 ;
        RECT 10.730 2174.490 11.910 2175.670 ;
        RECT 9.130 1996.090 10.310 1997.270 ;
        RECT 10.730 1996.090 11.910 1997.270 ;
        RECT 9.130 1994.490 10.310 1995.670 ;
        RECT 10.730 1994.490 11.910 1995.670 ;
        RECT 9.130 1816.090 10.310 1817.270 ;
        RECT 10.730 1816.090 11.910 1817.270 ;
        RECT 9.130 1814.490 10.310 1815.670 ;
        RECT 10.730 1814.490 11.910 1815.670 ;
        RECT 9.130 1636.090 10.310 1637.270 ;
        RECT 10.730 1636.090 11.910 1637.270 ;
        RECT 9.130 1634.490 10.310 1635.670 ;
        RECT 10.730 1634.490 11.910 1635.670 ;
        RECT 9.130 1456.090 10.310 1457.270 ;
        RECT 10.730 1456.090 11.910 1457.270 ;
        RECT 9.130 1454.490 10.310 1455.670 ;
        RECT 10.730 1454.490 11.910 1455.670 ;
        RECT 9.130 1276.090 10.310 1277.270 ;
        RECT 10.730 1276.090 11.910 1277.270 ;
        RECT 9.130 1274.490 10.310 1275.670 ;
        RECT 10.730 1274.490 11.910 1275.670 ;
        RECT 9.130 1096.090 10.310 1097.270 ;
        RECT 10.730 1096.090 11.910 1097.270 ;
        RECT 9.130 1094.490 10.310 1095.670 ;
        RECT 10.730 1094.490 11.910 1095.670 ;
        RECT 9.130 916.090 10.310 917.270 ;
        RECT 10.730 916.090 11.910 917.270 ;
        RECT 9.130 914.490 10.310 915.670 ;
        RECT 10.730 914.490 11.910 915.670 ;
        RECT 9.130 736.090 10.310 737.270 ;
        RECT 10.730 736.090 11.910 737.270 ;
        RECT 9.130 734.490 10.310 735.670 ;
        RECT 10.730 734.490 11.910 735.670 ;
        RECT 9.130 556.090 10.310 557.270 ;
        RECT 10.730 556.090 11.910 557.270 ;
        RECT 9.130 554.490 10.310 555.670 ;
        RECT 10.730 554.490 11.910 555.670 ;
        RECT 9.130 376.090 10.310 377.270 ;
        RECT 10.730 376.090 11.910 377.270 ;
        RECT 9.130 374.490 10.310 375.670 ;
        RECT 10.730 374.490 11.910 375.670 ;
        RECT 9.130 196.090 10.310 197.270 ;
        RECT 10.730 196.090 11.910 197.270 ;
        RECT 9.130 194.490 10.310 195.670 ;
        RECT 10.730 194.490 11.910 195.670 ;
        RECT 9.130 16.090 10.310 17.270 ;
        RECT 10.730 16.090 11.910 17.270 ;
        RECT 9.130 14.490 10.310 15.670 ;
        RECT 10.730 14.490 11.910 15.670 ;
        RECT 9.130 -4.460 10.310 -3.280 ;
        RECT 10.730 -4.460 11.910 -3.280 ;
        RECT 9.130 -6.060 10.310 -4.880 ;
        RECT 10.730 -6.060 11.910 -4.880 ;
        RECT 189.130 3524.560 190.310 3525.740 ;
        RECT 190.730 3524.560 191.910 3525.740 ;
        RECT 189.130 3522.960 190.310 3524.140 ;
        RECT 190.730 3522.960 191.910 3524.140 ;
        RECT 189.130 3436.090 190.310 3437.270 ;
        RECT 190.730 3436.090 191.910 3437.270 ;
        RECT 189.130 3434.490 190.310 3435.670 ;
        RECT 190.730 3434.490 191.910 3435.670 ;
        RECT 189.130 3256.090 190.310 3257.270 ;
        RECT 190.730 3256.090 191.910 3257.270 ;
        RECT 189.130 3254.490 190.310 3255.670 ;
        RECT 190.730 3254.490 191.910 3255.670 ;
        RECT 189.130 3076.090 190.310 3077.270 ;
        RECT 190.730 3076.090 191.910 3077.270 ;
        RECT 189.130 3074.490 190.310 3075.670 ;
        RECT 190.730 3074.490 191.910 3075.670 ;
        RECT 189.130 2896.090 190.310 2897.270 ;
        RECT 190.730 2896.090 191.910 2897.270 ;
        RECT 189.130 2894.490 190.310 2895.670 ;
        RECT 190.730 2894.490 191.910 2895.670 ;
        RECT 189.130 2716.090 190.310 2717.270 ;
        RECT 190.730 2716.090 191.910 2717.270 ;
        RECT 189.130 2714.490 190.310 2715.670 ;
        RECT 190.730 2714.490 191.910 2715.670 ;
        RECT 189.130 2536.090 190.310 2537.270 ;
        RECT 190.730 2536.090 191.910 2537.270 ;
        RECT 189.130 2534.490 190.310 2535.670 ;
        RECT 190.730 2534.490 191.910 2535.670 ;
        RECT 189.130 2356.090 190.310 2357.270 ;
        RECT 190.730 2356.090 191.910 2357.270 ;
        RECT 189.130 2354.490 190.310 2355.670 ;
        RECT 190.730 2354.490 191.910 2355.670 ;
        RECT 189.130 2176.090 190.310 2177.270 ;
        RECT 190.730 2176.090 191.910 2177.270 ;
        RECT 189.130 2174.490 190.310 2175.670 ;
        RECT 190.730 2174.490 191.910 2175.670 ;
        RECT 189.130 1996.090 190.310 1997.270 ;
        RECT 190.730 1996.090 191.910 1997.270 ;
        RECT 189.130 1994.490 190.310 1995.670 ;
        RECT 190.730 1994.490 191.910 1995.670 ;
        RECT 189.130 1816.090 190.310 1817.270 ;
        RECT 190.730 1816.090 191.910 1817.270 ;
        RECT 189.130 1814.490 190.310 1815.670 ;
        RECT 190.730 1814.490 191.910 1815.670 ;
        RECT 189.130 1636.090 190.310 1637.270 ;
        RECT 190.730 1636.090 191.910 1637.270 ;
        RECT 189.130 1634.490 190.310 1635.670 ;
        RECT 190.730 1634.490 191.910 1635.670 ;
        RECT 189.130 1456.090 190.310 1457.270 ;
        RECT 190.730 1456.090 191.910 1457.270 ;
        RECT 189.130 1454.490 190.310 1455.670 ;
        RECT 190.730 1454.490 191.910 1455.670 ;
        RECT 189.130 1276.090 190.310 1277.270 ;
        RECT 190.730 1276.090 191.910 1277.270 ;
        RECT 189.130 1274.490 190.310 1275.670 ;
        RECT 190.730 1274.490 191.910 1275.670 ;
        RECT 189.130 1096.090 190.310 1097.270 ;
        RECT 190.730 1096.090 191.910 1097.270 ;
        RECT 189.130 1094.490 190.310 1095.670 ;
        RECT 190.730 1094.490 191.910 1095.670 ;
        RECT 189.130 916.090 190.310 917.270 ;
        RECT 190.730 916.090 191.910 917.270 ;
        RECT 189.130 914.490 190.310 915.670 ;
        RECT 190.730 914.490 191.910 915.670 ;
        RECT 189.130 736.090 190.310 737.270 ;
        RECT 190.730 736.090 191.910 737.270 ;
        RECT 189.130 734.490 190.310 735.670 ;
        RECT 190.730 734.490 191.910 735.670 ;
        RECT 189.130 556.090 190.310 557.270 ;
        RECT 190.730 556.090 191.910 557.270 ;
        RECT 189.130 554.490 190.310 555.670 ;
        RECT 190.730 554.490 191.910 555.670 ;
        RECT 189.130 376.090 190.310 377.270 ;
        RECT 190.730 376.090 191.910 377.270 ;
        RECT 189.130 374.490 190.310 375.670 ;
        RECT 190.730 374.490 191.910 375.670 ;
        RECT 189.130 196.090 190.310 197.270 ;
        RECT 190.730 196.090 191.910 197.270 ;
        RECT 189.130 194.490 190.310 195.670 ;
        RECT 190.730 194.490 191.910 195.670 ;
        RECT 189.130 16.090 190.310 17.270 ;
        RECT 190.730 16.090 191.910 17.270 ;
        RECT 189.130 14.490 190.310 15.670 ;
        RECT 190.730 14.490 191.910 15.670 ;
        RECT 189.130 -4.460 190.310 -3.280 ;
        RECT 190.730 -4.460 191.910 -3.280 ;
        RECT 189.130 -6.060 190.310 -4.880 ;
        RECT 190.730 -6.060 191.910 -4.880 ;
        RECT 369.130 3524.560 370.310 3525.740 ;
        RECT 370.730 3524.560 371.910 3525.740 ;
        RECT 369.130 3522.960 370.310 3524.140 ;
        RECT 370.730 3522.960 371.910 3524.140 ;
        RECT 369.130 3436.090 370.310 3437.270 ;
        RECT 370.730 3436.090 371.910 3437.270 ;
        RECT 369.130 3434.490 370.310 3435.670 ;
        RECT 370.730 3434.490 371.910 3435.670 ;
        RECT 369.130 3256.090 370.310 3257.270 ;
        RECT 370.730 3256.090 371.910 3257.270 ;
        RECT 369.130 3254.490 370.310 3255.670 ;
        RECT 370.730 3254.490 371.910 3255.670 ;
        RECT 369.130 3076.090 370.310 3077.270 ;
        RECT 370.730 3076.090 371.910 3077.270 ;
        RECT 369.130 3074.490 370.310 3075.670 ;
        RECT 370.730 3074.490 371.910 3075.670 ;
        RECT 369.130 2896.090 370.310 2897.270 ;
        RECT 370.730 2896.090 371.910 2897.270 ;
        RECT 369.130 2894.490 370.310 2895.670 ;
        RECT 370.730 2894.490 371.910 2895.670 ;
        RECT 369.130 2716.090 370.310 2717.270 ;
        RECT 370.730 2716.090 371.910 2717.270 ;
        RECT 369.130 2714.490 370.310 2715.670 ;
        RECT 370.730 2714.490 371.910 2715.670 ;
        RECT 369.130 2536.090 370.310 2537.270 ;
        RECT 370.730 2536.090 371.910 2537.270 ;
        RECT 369.130 2534.490 370.310 2535.670 ;
        RECT 370.730 2534.490 371.910 2535.670 ;
        RECT 369.130 2356.090 370.310 2357.270 ;
        RECT 370.730 2356.090 371.910 2357.270 ;
        RECT 369.130 2354.490 370.310 2355.670 ;
        RECT 370.730 2354.490 371.910 2355.670 ;
        RECT 369.130 2176.090 370.310 2177.270 ;
        RECT 370.730 2176.090 371.910 2177.270 ;
        RECT 369.130 2174.490 370.310 2175.670 ;
        RECT 370.730 2174.490 371.910 2175.670 ;
        RECT 369.130 1996.090 370.310 1997.270 ;
        RECT 370.730 1996.090 371.910 1997.270 ;
        RECT 369.130 1994.490 370.310 1995.670 ;
        RECT 370.730 1994.490 371.910 1995.670 ;
        RECT 369.130 1816.090 370.310 1817.270 ;
        RECT 370.730 1816.090 371.910 1817.270 ;
        RECT 369.130 1814.490 370.310 1815.670 ;
        RECT 370.730 1814.490 371.910 1815.670 ;
        RECT 369.130 1636.090 370.310 1637.270 ;
        RECT 370.730 1636.090 371.910 1637.270 ;
        RECT 369.130 1634.490 370.310 1635.670 ;
        RECT 370.730 1634.490 371.910 1635.670 ;
        RECT 369.130 1456.090 370.310 1457.270 ;
        RECT 370.730 1456.090 371.910 1457.270 ;
        RECT 369.130 1454.490 370.310 1455.670 ;
        RECT 370.730 1454.490 371.910 1455.670 ;
        RECT 369.130 1276.090 370.310 1277.270 ;
        RECT 370.730 1276.090 371.910 1277.270 ;
        RECT 369.130 1274.490 370.310 1275.670 ;
        RECT 370.730 1274.490 371.910 1275.670 ;
        RECT 369.130 1096.090 370.310 1097.270 ;
        RECT 370.730 1096.090 371.910 1097.270 ;
        RECT 369.130 1094.490 370.310 1095.670 ;
        RECT 370.730 1094.490 371.910 1095.670 ;
        RECT 369.130 916.090 370.310 917.270 ;
        RECT 370.730 916.090 371.910 917.270 ;
        RECT 369.130 914.490 370.310 915.670 ;
        RECT 370.730 914.490 371.910 915.670 ;
        RECT 549.130 3524.560 550.310 3525.740 ;
        RECT 550.730 3524.560 551.910 3525.740 ;
        RECT 549.130 3522.960 550.310 3524.140 ;
        RECT 550.730 3522.960 551.910 3524.140 ;
        RECT 549.130 3436.090 550.310 3437.270 ;
        RECT 550.730 3436.090 551.910 3437.270 ;
        RECT 549.130 3434.490 550.310 3435.670 ;
        RECT 550.730 3434.490 551.910 3435.670 ;
        RECT 549.130 3256.090 550.310 3257.270 ;
        RECT 550.730 3256.090 551.910 3257.270 ;
        RECT 549.130 3254.490 550.310 3255.670 ;
        RECT 550.730 3254.490 551.910 3255.670 ;
        RECT 549.130 3076.090 550.310 3077.270 ;
        RECT 550.730 3076.090 551.910 3077.270 ;
        RECT 549.130 3074.490 550.310 3075.670 ;
        RECT 550.730 3074.490 551.910 3075.670 ;
        RECT 549.130 2896.090 550.310 2897.270 ;
        RECT 550.730 2896.090 551.910 2897.270 ;
        RECT 549.130 2894.490 550.310 2895.670 ;
        RECT 550.730 2894.490 551.910 2895.670 ;
        RECT 549.130 2716.090 550.310 2717.270 ;
        RECT 550.730 2716.090 551.910 2717.270 ;
        RECT 549.130 2714.490 550.310 2715.670 ;
        RECT 550.730 2714.490 551.910 2715.670 ;
        RECT 549.130 2536.090 550.310 2537.270 ;
        RECT 550.730 2536.090 551.910 2537.270 ;
        RECT 549.130 2534.490 550.310 2535.670 ;
        RECT 550.730 2534.490 551.910 2535.670 ;
        RECT 549.130 2356.090 550.310 2357.270 ;
        RECT 550.730 2356.090 551.910 2357.270 ;
        RECT 549.130 2354.490 550.310 2355.670 ;
        RECT 550.730 2354.490 551.910 2355.670 ;
        RECT 549.130 2176.090 550.310 2177.270 ;
        RECT 550.730 2176.090 551.910 2177.270 ;
        RECT 549.130 2174.490 550.310 2175.670 ;
        RECT 550.730 2174.490 551.910 2175.670 ;
        RECT 549.130 1996.090 550.310 1997.270 ;
        RECT 550.730 1996.090 551.910 1997.270 ;
        RECT 549.130 1994.490 550.310 1995.670 ;
        RECT 550.730 1994.490 551.910 1995.670 ;
        RECT 549.130 1816.090 550.310 1817.270 ;
        RECT 550.730 1816.090 551.910 1817.270 ;
        RECT 549.130 1814.490 550.310 1815.670 ;
        RECT 550.730 1814.490 551.910 1815.670 ;
        RECT 549.130 1636.090 550.310 1637.270 ;
        RECT 550.730 1636.090 551.910 1637.270 ;
        RECT 549.130 1634.490 550.310 1635.670 ;
        RECT 550.730 1634.490 551.910 1635.670 ;
        RECT 549.130 1456.090 550.310 1457.270 ;
        RECT 550.730 1456.090 551.910 1457.270 ;
        RECT 549.130 1454.490 550.310 1455.670 ;
        RECT 550.730 1454.490 551.910 1455.670 ;
        RECT 549.130 1276.090 550.310 1277.270 ;
        RECT 550.730 1276.090 551.910 1277.270 ;
        RECT 549.130 1274.490 550.310 1275.670 ;
        RECT 550.730 1274.490 551.910 1275.670 ;
        RECT 549.130 1096.090 550.310 1097.270 ;
        RECT 550.730 1096.090 551.910 1097.270 ;
        RECT 549.130 1094.490 550.310 1095.670 ;
        RECT 550.730 1094.490 551.910 1095.670 ;
        RECT 549.130 916.090 550.310 917.270 ;
        RECT 550.730 916.090 551.910 917.270 ;
        RECT 549.130 914.490 550.310 915.670 ;
        RECT 550.730 914.490 551.910 915.670 ;
        RECT 729.130 3524.560 730.310 3525.740 ;
        RECT 730.730 3524.560 731.910 3525.740 ;
        RECT 729.130 3522.960 730.310 3524.140 ;
        RECT 730.730 3522.960 731.910 3524.140 ;
        RECT 729.130 3436.090 730.310 3437.270 ;
        RECT 730.730 3436.090 731.910 3437.270 ;
        RECT 729.130 3434.490 730.310 3435.670 ;
        RECT 730.730 3434.490 731.910 3435.670 ;
        RECT 729.130 3256.090 730.310 3257.270 ;
        RECT 730.730 3256.090 731.910 3257.270 ;
        RECT 729.130 3254.490 730.310 3255.670 ;
        RECT 730.730 3254.490 731.910 3255.670 ;
        RECT 729.130 3076.090 730.310 3077.270 ;
        RECT 730.730 3076.090 731.910 3077.270 ;
        RECT 729.130 3074.490 730.310 3075.670 ;
        RECT 730.730 3074.490 731.910 3075.670 ;
        RECT 729.130 2896.090 730.310 2897.270 ;
        RECT 730.730 2896.090 731.910 2897.270 ;
        RECT 729.130 2894.490 730.310 2895.670 ;
        RECT 730.730 2894.490 731.910 2895.670 ;
        RECT 729.130 2716.090 730.310 2717.270 ;
        RECT 730.730 2716.090 731.910 2717.270 ;
        RECT 729.130 2714.490 730.310 2715.670 ;
        RECT 730.730 2714.490 731.910 2715.670 ;
        RECT 729.130 2536.090 730.310 2537.270 ;
        RECT 730.730 2536.090 731.910 2537.270 ;
        RECT 729.130 2534.490 730.310 2535.670 ;
        RECT 730.730 2534.490 731.910 2535.670 ;
        RECT 729.130 2356.090 730.310 2357.270 ;
        RECT 730.730 2356.090 731.910 2357.270 ;
        RECT 729.130 2354.490 730.310 2355.670 ;
        RECT 730.730 2354.490 731.910 2355.670 ;
        RECT 729.130 2176.090 730.310 2177.270 ;
        RECT 730.730 2176.090 731.910 2177.270 ;
        RECT 729.130 2174.490 730.310 2175.670 ;
        RECT 730.730 2174.490 731.910 2175.670 ;
        RECT 729.130 1996.090 730.310 1997.270 ;
        RECT 730.730 1996.090 731.910 1997.270 ;
        RECT 729.130 1994.490 730.310 1995.670 ;
        RECT 730.730 1994.490 731.910 1995.670 ;
        RECT 729.130 1816.090 730.310 1817.270 ;
        RECT 730.730 1816.090 731.910 1817.270 ;
        RECT 729.130 1814.490 730.310 1815.670 ;
        RECT 730.730 1814.490 731.910 1815.670 ;
        RECT 729.130 1636.090 730.310 1637.270 ;
        RECT 730.730 1636.090 731.910 1637.270 ;
        RECT 729.130 1634.490 730.310 1635.670 ;
        RECT 730.730 1634.490 731.910 1635.670 ;
        RECT 729.130 1456.090 730.310 1457.270 ;
        RECT 730.730 1456.090 731.910 1457.270 ;
        RECT 729.130 1454.490 730.310 1455.670 ;
        RECT 730.730 1454.490 731.910 1455.670 ;
        RECT 729.130 1276.090 730.310 1277.270 ;
        RECT 730.730 1276.090 731.910 1277.270 ;
        RECT 729.130 1274.490 730.310 1275.670 ;
        RECT 730.730 1274.490 731.910 1275.670 ;
        RECT 729.130 1096.090 730.310 1097.270 ;
        RECT 730.730 1096.090 731.910 1097.270 ;
        RECT 729.130 1094.490 730.310 1095.670 ;
        RECT 730.730 1094.490 731.910 1095.670 ;
        RECT 729.130 916.090 730.310 917.270 ;
        RECT 730.730 916.090 731.910 917.270 ;
        RECT 729.130 914.490 730.310 915.670 ;
        RECT 730.730 914.490 731.910 915.670 ;
        RECT 369.130 736.090 370.310 737.270 ;
        RECT 370.730 736.090 371.910 737.270 ;
        RECT 369.130 734.490 370.310 735.670 ;
        RECT 370.730 734.490 371.910 735.670 ;
        RECT 369.130 556.090 370.310 557.270 ;
        RECT 370.730 556.090 371.910 557.270 ;
        RECT 369.130 554.490 370.310 555.670 ;
        RECT 370.730 554.490 371.910 555.670 ;
        RECT 421.250 735.015 422.430 736.195 ;
        RECT 421.250 556.090 422.430 557.270 ;
        RECT 421.250 554.490 422.430 555.670 ;
        RECT 574.850 735.015 576.030 736.195 ;
        RECT 574.850 556.090 576.030 557.270 ;
        RECT 574.850 554.490 576.030 555.670 ;
        RECT 729.130 736.090 730.310 737.270 ;
        RECT 730.730 736.090 731.910 737.270 ;
        RECT 729.130 734.490 730.310 735.670 ;
        RECT 730.730 734.490 731.910 735.670 ;
        RECT 729.130 556.090 730.310 557.270 ;
        RECT 730.730 556.090 731.910 557.270 ;
        RECT 729.130 554.490 730.310 555.670 ;
        RECT 730.730 554.490 731.910 555.670 ;
        RECT 369.130 376.090 370.310 377.270 ;
        RECT 370.730 376.090 371.910 377.270 ;
        RECT 369.130 374.490 370.310 375.670 ;
        RECT 370.730 374.490 371.910 375.670 ;
        RECT 369.130 196.090 370.310 197.270 ;
        RECT 370.730 196.090 371.910 197.270 ;
        RECT 369.130 194.490 370.310 195.670 ;
        RECT 370.730 194.490 371.910 195.670 ;
        RECT 369.130 16.090 370.310 17.270 ;
        RECT 370.730 16.090 371.910 17.270 ;
        RECT 369.130 14.490 370.310 15.670 ;
        RECT 370.730 14.490 371.910 15.670 ;
        RECT 369.130 -4.460 370.310 -3.280 ;
        RECT 370.730 -4.460 371.910 -3.280 ;
        RECT 369.130 -6.060 370.310 -4.880 ;
        RECT 370.730 -6.060 371.910 -4.880 ;
        RECT 549.130 376.090 550.310 377.270 ;
        RECT 550.730 376.090 551.910 377.270 ;
        RECT 549.130 374.490 550.310 375.670 ;
        RECT 550.730 374.490 551.910 375.670 ;
        RECT 549.130 196.090 550.310 197.270 ;
        RECT 550.730 196.090 551.910 197.270 ;
        RECT 549.130 194.490 550.310 195.670 ;
        RECT 550.730 194.490 551.910 195.670 ;
        RECT 549.130 16.090 550.310 17.270 ;
        RECT 550.730 16.090 551.910 17.270 ;
        RECT 549.130 14.490 550.310 15.670 ;
        RECT 550.730 14.490 551.910 15.670 ;
        RECT 549.130 -4.460 550.310 -3.280 ;
        RECT 550.730 -4.460 551.910 -3.280 ;
        RECT 549.130 -6.060 550.310 -4.880 ;
        RECT 550.730 -6.060 551.910 -4.880 ;
        RECT 729.130 376.090 730.310 377.270 ;
        RECT 730.730 376.090 731.910 377.270 ;
        RECT 729.130 374.490 730.310 375.670 ;
        RECT 730.730 374.490 731.910 375.670 ;
        RECT 729.130 196.090 730.310 197.270 ;
        RECT 730.730 196.090 731.910 197.270 ;
        RECT 729.130 194.490 730.310 195.670 ;
        RECT 730.730 194.490 731.910 195.670 ;
        RECT 729.130 16.090 730.310 17.270 ;
        RECT 730.730 16.090 731.910 17.270 ;
        RECT 729.130 14.490 730.310 15.670 ;
        RECT 730.730 14.490 731.910 15.670 ;
        RECT 729.130 -4.460 730.310 -3.280 ;
        RECT 730.730 -4.460 731.910 -3.280 ;
        RECT 729.130 -6.060 730.310 -4.880 ;
        RECT 730.730 -6.060 731.910 -4.880 ;
        RECT 909.130 3524.560 910.310 3525.740 ;
        RECT 910.730 3524.560 911.910 3525.740 ;
        RECT 909.130 3522.960 910.310 3524.140 ;
        RECT 910.730 3522.960 911.910 3524.140 ;
        RECT 909.130 3436.090 910.310 3437.270 ;
        RECT 910.730 3436.090 911.910 3437.270 ;
        RECT 909.130 3434.490 910.310 3435.670 ;
        RECT 910.730 3434.490 911.910 3435.670 ;
        RECT 909.130 3256.090 910.310 3257.270 ;
        RECT 910.730 3256.090 911.910 3257.270 ;
        RECT 909.130 3254.490 910.310 3255.670 ;
        RECT 910.730 3254.490 911.910 3255.670 ;
        RECT 909.130 3076.090 910.310 3077.270 ;
        RECT 910.730 3076.090 911.910 3077.270 ;
        RECT 909.130 3074.490 910.310 3075.670 ;
        RECT 910.730 3074.490 911.910 3075.670 ;
        RECT 909.130 2896.090 910.310 2897.270 ;
        RECT 910.730 2896.090 911.910 2897.270 ;
        RECT 909.130 2894.490 910.310 2895.670 ;
        RECT 910.730 2894.490 911.910 2895.670 ;
        RECT 909.130 2716.090 910.310 2717.270 ;
        RECT 910.730 2716.090 911.910 2717.270 ;
        RECT 909.130 2714.490 910.310 2715.670 ;
        RECT 910.730 2714.490 911.910 2715.670 ;
        RECT 909.130 2536.090 910.310 2537.270 ;
        RECT 910.730 2536.090 911.910 2537.270 ;
        RECT 909.130 2534.490 910.310 2535.670 ;
        RECT 910.730 2534.490 911.910 2535.670 ;
        RECT 909.130 2356.090 910.310 2357.270 ;
        RECT 910.730 2356.090 911.910 2357.270 ;
        RECT 909.130 2354.490 910.310 2355.670 ;
        RECT 910.730 2354.490 911.910 2355.670 ;
        RECT 909.130 2176.090 910.310 2177.270 ;
        RECT 910.730 2176.090 911.910 2177.270 ;
        RECT 909.130 2174.490 910.310 2175.670 ;
        RECT 910.730 2174.490 911.910 2175.670 ;
        RECT 909.130 1996.090 910.310 1997.270 ;
        RECT 910.730 1996.090 911.910 1997.270 ;
        RECT 909.130 1994.490 910.310 1995.670 ;
        RECT 910.730 1994.490 911.910 1995.670 ;
        RECT 909.130 1816.090 910.310 1817.270 ;
        RECT 910.730 1816.090 911.910 1817.270 ;
        RECT 909.130 1814.490 910.310 1815.670 ;
        RECT 910.730 1814.490 911.910 1815.670 ;
        RECT 909.130 1636.090 910.310 1637.270 ;
        RECT 910.730 1636.090 911.910 1637.270 ;
        RECT 909.130 1634.490 910.310 1635.670 ;
        RECT 910.730 1634.490 911.910 1635.670 ;
        RECT 909.130 1456.090 910.310 1457.270 ;
        RECT 910.730 1456.090 911.910 1457.270 ;
        RECT 909.130 1454.490 910.310 1455.670 ;
        RECT 910.730 1454.490 911.910 1455.670 ;
        RECT 909.130 1276.090 910.310 1277.270 ;
        RECT 910.730 1276.090 911.910 1277.270 ;
        RECT 909.130 1274.490 910.310 1275.670 ;
        RECT 910.730 1274.490 911.910 1275.670 ;
        RECT 909.130 1096.090 910.310 1097.270 ;
        RECT 910.730 1096.090 911.910 1097.270 ;
        RECT 909.130 1094.490 910.310 1095.670 ;
        RECT 910.730 1094.490 911.910 1095.670 ;
        RECT 909.130 916.090 910.310 917.270 ;
        RECT 910.730 916.090 911.910 917.270 ;
        RECT 909.130 914.490 910.310 915.670 ;
        RECT 910.730 914.490 911.910 915.670 ;
        RECT 909.130 736.090 910.310 737.270 ;
        RECT 910.730 736.090 911.910 737.270 ;
        RECT 909.130 734.490 910.310 735.670 ;
        RECT 910.730 734.490 911.910 735.670 ;
        RECT 909.130 556.090 910.310 557.270 ;
        RECT 910.730 556.090 911.910 557.270 ;
        RECT 909.130 554.490 910.310 555.670 ;
        RECT 910.730 554.490 911.910 555.670 ;
        RECT 909.130 376.090 910.310 377.270 ;
        RECT 910.730 376.090 911.910 377.270 ;
        RECT 909.130 374.490 910.310 375.670 ;
        RECT 910.730 374.490 911.910 375.670 ;
        RECT 909.130 196.090 910.310 197.270 ;
        RECT 910.730 196.090 911.910 197.270 ;
        RECT 909.130 194.490 910.310 195.670 ;
        RECT 910.730 194.490 911.910 195.670 ;
        RECT 909.130 16.090 910.310 17.270 ;
        RECT 910.730 16.090 911.910 17.270 ;
        RECT 909.130 14.490 910.310 15.670 ;
        RECT 910.730 14.490 911.910 15.670 ;
        RECT 909.130 -4.460 910.310 -3.280 ;
        RECT 910.730 -4.460 911.910 -3.280 ;
        RECT 909.130 -6.060 910.310 -4.880 ;
        RECT 910.730 -6.060 911.910 -4.880 ;
        RECT 1089.130 3524.560 1090.310 3525.740 ;
        RECT 1090.730 3524.560 1091.910 3525.740 ;
        RECT 1089.130 3522.960 1090.310 3524.140 ;
        RECT 1090.730 3522.960 1091.910 3524.140 ;
        RECT 1089.130 3436.090 1090.310 3437.270 ;
        RECT 1090.730 3436.090 1091.910 3437.270 ;
        RECT 1089.130 3434.490 1090.310 3435.670 ;
        RECT 1090.730 3434.490 1091.910 3435.670 ;
        RECT 1089.130 3256.090 1090.310 3257.270 ;
        RECT 1090.730 3256.090 1091.910 3257.270 ;
        RECT 1089.130 3254.490 1090.310 3255.670 ;
        RECT 1090.730 3254.490 1091.910 3255.670 ;
        RECT 1089.130 3076.090 1090.310 3077.270 ;
        RECT 1090.730 3076.090 1091.910 3077.270 ;
        RECT 1089.130 3074.490 1090.310 3075.670 ;
        RECT 1090.730 3074.490 1091.910 3075.670 ;
        RECT 1089.130 2896.090 1090.310 2897.270 ;
        RECT 1090.730 2896.090 1091.910 2897.270 ;
        RECT 1089.130 2894.490 1090.310 2895.670 ;
        RECT 1090.730 2894.490 1091.910 2895.670 ;
        RECT 1089.130 2716.090 1090.310 2717.270 ;
        RECT 1090.730 2716.090 1091.910 2717.270 ;
        RECT 1089.130 2714.490 1090.310 2715.670 ;
        RECT 1090.730 2714.490 1091.910 2715.670 ;
        RECT 1089.130 2536.090 1090.310 2537.270 ;
        RECT 1090.730 2536.090 1091.910 2537.270 ;
        RECT 1089.130 2534.490 1090.310 2535.670 ;
        RECT 1090.730 2534.490 1091.910 2535.670 ;
        RECT 1089.130 2356.090 1090.310 2357.270 ;
        RECT 1090.730 2356.090 1091.910 2357.270 ;
        RECT 1089.130 2354.490 1090.310 2355.670 ;
        RECT 1090.730 2354.490 1091.910 2355.670 ;
        RECT 1089.130 2176.090 1090.310 2177.270 ;
        RECT 1090.730 2176.090 1091.910 2177.270 ;
        RECT 1089.130 2174.490 1090.310 2175.670 ;
        RECT 1090.730 2174.490 1091.910 2175.670 ;
        RECT 1089.130 1996.090 1090.310 1997.270 ;
        RECT 1090.730 1996.090 1091.910 1997.270 ;
        RECT 1089.130 1994.490 1090.310 1995.670 ;
        RECT 1090.730 1994.490 1091.910 1995.670 ;
        RECT 1089.130 1816.090 1090.310 1817.270 ;
        RECT 1090.730 1816.090 1091.910 1817.270 ;
        RECT 1089.130 1814.490 1090.310 1815.670 ;
        RECT 1090.730 1814.490 1091.910 1815.670 ;
        RECT 1089.130 1636.090 1090.310 1637.270 ;
        RECT 1090.730 1636.090 1091.910 1637.270 ;
        RECT 1089.130 1634.490 1090.310 1635.670 ;
        RECT 1090.730 1634.490 1091.910 1635.670 ;
        RECT 1089.130 1456.090 1090.310 1457.270 ;
        RECT 1090.730 1456.090 1091.910 1457.270 ;
        RECT 1089.130 1454.490 1090.310 1455.670 ;
        RECT 1090.730 1454.490 1091.910 1455.670 ;
        RECT 1089.130 1276.090 1090.310 1277.270 ;
        RECT 1090.730 1276.090 1091.910 1277.270 ;
        RECT 1089.130 1274.490 1090.310 1275.670 ;
        RECT 1090.730 1274.490 1091.910 1275.670 ;
        RECT 1089.130 1096.090 1090.310 1097.270 ;
        RECT 1090.730 1096.090 1091.910 1097.270 ;
        RECT 1089.130 1094.490 1090.310 1095.670 ;
        RECT 1090.730 1094.490 1091.910 1095.670 ;
        RECT 1089.130 916.090 1090.310 917.270 ;
        RECT 1090.730 916.090 1091.910 917.270 ;
        RECT 1089.130 914.490 1090.310 915.670 ;
        RECT 1090.730 914.490 1091.910 915.670 ;
        RECT 1089.130 736.090 1090.310 737.270 ;
        RECT 1090.730 736.090 1091.910 737.270 ;
        RECT 1089.130 734.490 1090.310 735.670 ;
        RECT 1090.730 734.490 1091.910 735.670 ;
        RECT 1089.130 556.090 1090.310 557.270 ;
        RECT 1090.730 556.090 1091.910 557.270 ;
        RECT 1089.130 554.490 1090.310 555.670 ;
        RECT 1090.730 554.490 1091.910 555.670 ;
        RECT 1089.130 376.090 1090.310 377.270 ;
        RECT 1090.730 376.090 1091.910 377.270 ;
        RECT 1089.130 374.490 1090.310 375.670 ;
        RECT 1090.730 374.490 1091.910 375.670 ;
        RECT 1089.130 196.090 1090.310 197.270 ;
        RECT 1090.730 196.090 1091.910 197.270 ;
        RECT 1089.130 194.490 1090.310 195.670 ;
        RECT 1090.730 194.490 1091.910 195.670 ;
        RECT 1089.130 16.090 1090.310 17.270 ;
        RECT 1090.730 16.090 1091.910 17.270 ;
        RECT 1089.130 14.490 1090.310 15.670 ;
        RECT 1090.730 14.490 1091.910 15.670 ;
        RECT 1089.130 -4.460 1090.310 -3.280 ;
        RECT 1090.730 -4.460 1091.910 -3.280 ;
        RECT 1089.130 -6.060 1090.310 -4.880 ;
        RECT 1090.730 -6.060 1091.910 -4.880 ;
        RECT 1269.130 3524.560 1270.310 3525.740 ;
        RECT 1270.730 3524.560 1271.910 3525.740 ;
        RECT 1269.130 3522.960 1270.310 3524.140 ;
        RECT 1270.730 3522.960 1271.910 3524.140 ;
        RECT 1269.130 3436.090 1270.310 3437.270 ;
        RECT 1270.730 3436.090 1271.910 3437.270 ;
        RECT 1269.130 3434.490 1270.310 3435.670 ;
        RECT 1270.730 3434.490 1271.910 3435.670 ;
        RECT 1269.130 3256.090 1270.310 3257.270 ;
        RECT 1270.730 3256.090 1271.910 3257.270 ;
        RECT 1269.130 3254.490 1270.310 3255.670 ;
        RECT 1270.730 3254.490 1271.910 3255.670 ;
        RECT 1269.130 3076.090 1270.310 3077.270 ;
        RECT 1270.730 3076.090 1271.910 3077.270 ;
        RECT 1269.130 3074.490 1270.310 3075.670 ;
        RECT 1270.730 3074.490 1271.910 3075.670 ;
        RECT 1269.130 2896.090 1270.310 2897.270 ;
        RECT 1270.730 2896.090 1271.910 2897.270 ;
        RECT 1269.130 2894.490 1270.310 2895.670 ;
        RECT 1270.730 2894.490 1271.910 2895.670 ;
        RECT 1269.130 2716.090 1270.310 2717.270 ;
        RECT 1270.730 2716.090 1271.910 2717.270 ;
        RECT 1269.130 2714.490 1270.310 2715.670 ;
        RECT 1270.730 2714.490 1271.910 2715.670 ;
        RECT 1269.130 2536.090 1270.310 2537.270 ;
        RECT 1270.730 2536.090 1271.910 2537.270 ;
        RECT 1269.130 2534.490 1270.310 2535.670 ;
        RECT 1270.730 2534.490 1271.910 2535.670 ;
        RECT 1269.130 2356.090 1270.310 2357.270 ;
        RECT 1270.730 2356.090 1271.910 2357.270 ;
        RECT 1269.130 2354.490 1270.310 2355.670 ;
        RECT 1270.730 2354.490 1271.910 2355.670 ;
        RECT 1269.130 2176.090 1270.310 2177.270 ;
        RECT 1270.730 2176.090 1271.910 2177.270 ;
        RECT 1269.130 2174.490 1270.310 2175.670 ;
        RECT 1270.730 2174.490 1271.910 2175.670 ;
        RECT 1269.130 1996.090 1270.310 1997.270 ;
        RECT 1270.730 1996.090 1271.910 1997.270 ;
        RECT 1269.130 1994.490 1270.310 1995.670 ;
        RECT 1270.730 1994.490 1271.910 1995.670 ;
        RECT 1269.130 1816.090 1270.310 1817.270 ;
        RECT 1270.730 1816.090 1271.910 1817.270 ;
        RECT 1269.130 1814.490 1270.310 1815.670 ;
        RECT 1270.730 1814.490 1271.910 1815.670 ;
        RECT 1269.130 1636.090 1270.310 1637.270 ;
        RECT 1270.730 1636.090 1271.910 1637.270 ;
        RECT 1269.130 1634.490 1270.310 1635.670 ;
        RECT 1270.730 1634.490 1271.910 1635.670 ;
        RECT 1269.130 1456.090 1270.310 1457.270 ;
        RECT 1270.730 1456.090 1271.910 1457.270 ;
        RECT 1269.130 1454.490 1270.310 1455.670 ;
        RECT 1270.730 1454.490 1271.910 1455.670 ;
        RECT 1269.130 1276.090 1270.310 1277.270 ;
        RECT 1270.730 1276.090 1271.910 1277.270 ;
        RECT 1269.130 1274.490 1270.310 1275.670 ;
        RECT 1270.730 1274.490 1271.910 1275.670 ;
        RECT 1269.130 1096.090 1270.310 1097.270 ;
        RECT 1270.730 1096.090 1271.910 1097.270 ;
        RECT 1269.130 1094.490 1270.310 1095.670 ;
        RECT 1270.730 1094.490 1271.910 1095.670 ;
        RECT 1269.130 916.090 1270.310 917.270 ;
        RECT 1270.730 916.090 1271.910 917.270 ;
        RECT 1269.130 914.490 1270.310 915.670 ;
        RECT 1270.730 914.490 1271.910 915.670 ;
        RECT 1269.130 736.090 1270.310 737.270 ;
        RECT 1270.730 736.090 1271.910 737.270 ;
        RECT 1269.130 734.490 1270.310 735.670 ;
        RECT 1270.730 734.490 1271.910 735.670 ;
        RECT 1269.130 556.090 1270.310 557.270 ;
        RECT 1270.730 556.090 1271.910 557.270 ;
        RECT 1269.130 554.490 1270.310 555.670 ;
        RECT 1270.730 554.490 1271.910 555.670 ;
        RECT 1269.130 376.090 1270.310 377.270 ;
        RECT 1270.730 376.090 1271.910 377.270 ;
        RECT 1269.130 374.490 1270.310 375.670 ;
        RECT 1270.730 374.490 1271.910 375.670 ;
        RECT 1269.130 196.090 1270.310 197.270 ;
        RECT 1270.730 196.090 1271.910 197.270 ;
        RECT 1269.130 194.490 1270.310 195.670 ;
        RECT 1270.730 194.490 1271.910 195.670 ;
        RECT 1269.130 16.090 1270.310 17.270 ;
        RECT 1270.730 16.090 1271.910 17.270 ;
        RECT 1269.130 14.490 1270.310 15.670 ;
        RECT 1270.730 14.490 1271.910 15.670 ;
        RECT 1269.130 -4.460 1270.310 -3.280 ;
        RECT 1270.730 -4.460 1271.910 -3.280 ;
        RECT 1269.130 -6.060 1270.310 -4.880 ;
        RECT 1270.730 -6.060 1271.910 -4.880 ;
        RECT 1449.130 3524.560 1450.310 3525.740 ;
        RECT 1450.730 3524.560 1451.910 3525.740 ;
        RECT 1449.130 3522.960 1450.310 3524.140 ;
        RECT 1450.730 3522.960 1451.910 3524.140 ;
        RECT 1449.130 3436.090 1450.310 3437.270 ;
        RECT 1450.730 3436.090 1451.910 3437.270 ;
        RECT 1449.130 3434.490 1450.310 3435.670 ;
        RECT 1450.730 3434.490 1451.910 3435.670 ;
        RECT 1449.130 3256.090 1450.310 3257.270 ;
        RECT 1450.730 3256.090 1451.910 3257.270 ;
        RECT 1449.130 3254.490 1450.310 3255.670 ;
        RECT 1450.730 3254.490 1451.910 3255.670 ;
        RECT 1449.130 3076.090 1450.310 3077.270 ;
        RECT 1450.730 3076.090 1451.910 3077.270 ;
        RECT 1449.130 3074.490 1450.310 3075.670 ;
        RECT 1450.730 3074.490 1451.910 3075.670 ;
        RECT 1449.130 2896.090 1450.310 2897.270 ;
        RECT 1450.730 2896.090 1451.910 2897.270 ;
        RECT 1449.130 2894.490 1450.310 2895.670 ;
        RECT 1450.730 2894.490 1451.910 2895.670 ;
        RECT 1449.130 2716.090 1450.310 2717.270 ;
        RECT 1450.730 2716.090 1451.910 2717.270 ;
        RECT 1449.130 2714.490 1450.310 2715.670 ;
        RECT 1450.730 2714.490 1451.910 2715.670 ;
        RECT 1449.130 2536.090 1450.310 2537.270 ;
        RECT 1450.730 2536.090 1451.910 2537.270 ;
        RECT 1449.130 2534.490 1450.310 2535.670 ;
        RECT 1450.730 2534.490 1451.910 2535.670 ;
        RECT 1449.130 2356.090 1450.310 2357.270 ;
        RECT 1450.730 2356.090 1451.910 2357.270 ;
        RECT 1449.130 2354.490 1450.310 2355.670 ;
        RECT 1450.730 2354.490 1451.910 2355.670 ;
        RECT 1449.130 2176.090 1450.310 2177.270 ;
        RECT 1450.730 2176.090 1451.910 2177.270 ;
        RECT 1449.130 2174.490 1450.310 2175.670 ;
        RECT 1450.730 2174.490 1451.910 2175.670 ;
        RECT 1449.130 1996.090 1450.310 1997.270 ;
        RECT 1450.730 1996.090 1451.910 1997.270 ;
        RECT 1449.130 1994.490 1450.310 1995.670 ;
        RECT 1450.730 1994.490 1451.910 1995.670 ;
        RECT 1449.130 1816.090 1450.310 1817.270 ;
        RECT 1450.730 1816.090 1451.910 1817.270 ;
        RECT 1449.130 1814.490 1450.310 1815.670 ;
        RECT 1450.730 1814.490 1451.910 1815.670 ;
        RECT 1449.130 1636.090 1450.310 1637.270 ;
        RECT 1450.730 1636.090 1451.910 1637.270 ;
        RECT 1449.130 1634.490 1450.310 1635.670 ;
        RECT 1450.730 1634.490 1451.910 1635.670 ;
        RECT 1449.130 1456.090 1450.310 1457.270 ;
        RECT 1450.730 1456.090 1451.910 1457.270 ;
        RECT 1449.130 1454.490 1450.310 1455.670 ;
        RECT 1450.730 1454.490 1451.910 1455.670 ;
        RECT 1449.130 1276.090 1450.310 1277.270 ;
        RECT 1450.730 1276.090 1451.910 1277.270 ;
        RECT 1449.130 1274.490 1450.310 1275.670 ;
        RECT 1450.730 1274.490 1451.910 1275.670 ;
        RECT 1449.130 1096.090 1450.310 1097.270 ;
        RECT 1450.730 1096.090 1451.910 1097.270 ;
        RECT 1449.130 1094.490 1450.310 1095.670 ;
        RECT 1450.730 1094.490 1451.910 1095.670 ;
        RECT 1449.130 916.090 1450.310 917.270 ;
        RECT 1450.730 916.090 1451.910 917.270 ;
        RECT 1449.130 914.490 1450.310 915.670 ;
        RECT 1450.730 914.490 1451.910 915.670 ;
        RECT 1449.130 736.090 1450.310 737.270 ;
        RECT 1450.730 736.090 1451.910 737.270 ;
        RECT 1449.130 734.490 1450.310 735.670 ;
        RECT 1450.730 734.490 1451.910 735.670 ;
        RECT 1449.130 556.090 1450.310 557.270 ;
        RECT 1450.730 556.090 1451.910 557.270 ;
        RECT 1449.130 554.490 1450.310 555.670 ;
        RECT 1450.730 554.490 1451.910 555.670 ;
        RECT 1449.130 376.090 1450.310 377.270 ;
        RECT 1450.730 376.090 1451.910 377.270 ;
        RECT 1449.130 374.490 1450.310 375.670 ;
        RECT 1450.730 374.490 1451.910 375.670 ;
        RECT 1449.130 196.090 1450.310 197.270 ;
        RECT 1450.730 196.090 1451.910 197.270 ;
        RECT 1449.130 194.490 1450.310 195.670 ;
        RECT 1450.730 194.490 1451.910 195.670 ;
        RECT 1449.130 16.090 1450.310 17.270 ;
        RECT 1450.730 16.090 1451.910 17.270 ;
        RECT 1449.130 14.490 1450.310 15.670 ;
        RECT 1450.730 14.490 1451.910 15.670 ;
        RECT 1449.130 -4.460 1450.310 -3.280 ;
        RECT 1450.730 -4.460 1451.910 -3.280 ;
        RECT 1449.130 -6.060 1450.310 -4.880 ;
        RECT 1450.730 -6.060 1451.910 -4.880 ;
        RECT 1629.130 3524.560 1630.310 3525.740 ;
        RECT 1630.730 3524.560 1631.910 3525.740 ;
        RECT 1629.130 3522.960 1630.310 3524.140 ;
        RECT 1630.730 3522.960 1631.910 3524.140 ;
        RECT 1629.130 3436.090 1630.310 3437.270 ;
        RECT 1630.730 3436.090 1631.910 3437.270 ;
        RECT 1629.130 3434.490 1630.310 3435.670 ;
        RECT 1630.730 3434.490 1631.910 3435.670 ;
        RECT 1629.130 3256.090 1630.310 3257.270 ;
        RECT 1630.730 3256.090 1631.910 3257.270 ;
        RECT 1629.130 3254.490 1630.310 3255.670 ;
        RECT 1630.730 3254.490 1631.910 3255.670 ;
        RECT 1629.130 3076.090 1630.310 3077.270 ;
        RECT 1630.730 3076.090 1631.910 3077.270 ;
        RECT 1629.130 3074.490 1630.310 3075.670 ;
        RECT 1630.730 3074.490 1631.910 3075.670 ;
        RECT 1629.130 2896.090 1630.310 2897.270 ;
        RECT 1630.730 2896.090 1631.910 2897.270 ;
        RECT 1629.130 2894.490 1630.310 2895.670 ;
        RECT 1630.730 2894.490 1631.910 2895.670 ;
        RECT 1629.130 2716.090 1630.310 2717.270 ;
        RECT 1630.730 2716.090 1631.910 2717.270 ;
        RECT 1629.130 2714.490 1630.310 2715.670 ;
        RECT 1630.730 2714.490 1631.910 2715.670 ;
        RECT 1629.130 2536.090 1630.310 2537.270 ;
        RECT 1630.730 2536.090 1631.910 2537.270 ;
        RECT 1629.130 2534.490 1630.310 2535.670 ;
        RECT 1630.730 2534.490 1631.910 2535.670 ;
        RECT 1629.130 2356.090 1630.310 2357.270 ;
        RECT 1630.730 2356.090 1631.910 2357.270 ;
        RECT 1629.130 2354.490 1630.310 2355.670 ;
        RECT 1630.730 2354.490 1631.910 2355.670 ;
        RECT 1629.130 2176.090 1630.310 2177.270 ;
        RECT 1630.730 2176.090 1631.910 2177.270 ;
        RECT 1629.130 2174.490 1630.310 2175.670 ;
        RECT 1630.730 2174.490 1631.910 2175.670 ;
        RECT 1629.130 1996.090 1630.310 1997.270 ;
        RECT 1630.730 1996.090 1631.910 1997.270 ;
        RECT 1629.130 1994.490 1630.310 1995.670 ;
        RECT 1630.730 1994.490 1631.910 1995.670 ;
        RECT 1629.130 1816.090 1630.310 1817.270 ;
        RECT 1630.730 1816.090 1631.910 1817.270 ;
        RECT 1629.130 1814.490 1630.310 1815.670 ;
        RECT 1630.730 1814.490 1631.910 1815.670 ;
        RECT 1629.130 1636.090 1630.310 1637.270 ;
        RECT 1630.730 1636.090 1631.910 1637.270 ;
        RECT 1629.130 1634.490 1630.310 1635.670 ;
        RECT 1630.730 1634.490 1631.910 1635.670 ;
        RECT 1629.130 1456.090 1630.310 1457.270 ;
        RECT 1630.730 1456.090 1631.910 1457.270 ;
        RECT 1629.130 1454.490 1630.310 1455.670 ;
        RECT 1630.730 1454.490 1631.910 1455.670 ;
        RECT 1629.130 1276.090 1630.310 1277.270 ;
        RECT 1630.730 1276.090 1631.910 1277.270 ;
        RECT 1629.130 1274.490 1630.310 1275.670 ;
        RECT 1630.730 1274.490 1631.910 1275.670 ;
        RECT 1629.130 1096.090 1630.310 1097.270 ;
        RECT 1630.730 1096.090 1631.910 1097.270 ;
        RECT 1629.130 1094.490 1630.310 1095.670 ;
        RECT 1630.730 1094.490 1631.910 1095.670 ;
        RECT 1629.130 916.090 1630.310 917.270 ;
        RECT 1630.730 916.090 1631.910 917.270 ;
        RECT 1629.130 914.490 1630.310 915.670 ;
        RECT 1630.730 914.490 1631.910 915.670 ;
        RECT 1629.130 736.090 1630.310 737.270 ;
        RECT 1630.730 736.090 1631.910 737.270 ;
        RECT 1629.130 734.490 1630.310 735.670 ;
        RECT 1630.730 734.490 1631.910 735.670 ;
        RECT 1629.130 556.090 1630.310 557.270 ;
        RECT 1630.730 556.090 1631.910 557.270 ;
        RECT 1629.130 554.490 1630.310 555.670 ;
        RECT 1630.730 554.490 1631.910 555.670 ;
        RECT 1629.130 376.090 1630.310 377.270 ;
        RECT 1630.730 376.090 1631.910 377.270 ;
        RECT 1629.130 374.490 1630.310 375.670 ;
        RECT 1630.730 374.490 1631.910 375.670 ;
        RECT 1629.130 196.090 1630.310 197.270 ;
        RECT 1630.730 196.090 1631.910 197.270 ;
        RECT 1629.130 194.490 1630.310 195.670 ;
        RECT 1630.730 194.490 1631.910 195.670 ;
        RECT 1629.130 16.090 1630.310 17.270 ;
        RECT 1630.730 16.090 1631.910 17.270 ;
        RECT 1629.130 14.490 1630.310 15.670 ;
        RECT 1630.730 14.490 1631.910 15.670 ;
        RECT 1629.130 -4.460 1630.310 -3.280 ;
        RECT 1630.730 -4.460 1631.910 -3.280 ;
        RECT 1629.130 -6.060 1630.310 -4.880 ;
        RECT 1630.730 -6.060 1631.910 -4.880 ;
        RECT 1809.130 3524.560 1810.310 3525.740 ;
        RECT 1810.730 3524.560 1811.910 3525.740 ;
        RECT 1809.130 3522.960 1810.310 3524.140 ;
        RECT 1810.730 3522.960 1811.910 3524.140 ;
        RECT 1809.130 3436.090 1810.310 3437.270 ;
        RECT 1810.730 3436.090 1811.910 3437.270 ;
        RECT 1809.130 3434.490 1810.310 3435.670 ;
        RECT 1810.730 3434.490 1811.910 3435.670 ;
        RECT 1809.130 3256.090 1810.310 3257.270 ;
        RECT 1810.730 3256.090 1811.910 3257.270 ;
        RECT 1809.130 3254.490 1810.310 3255.670 ;
        RECT 1810.730 3254.490 1811.910 3255.670 ;
        RECT 1809.130 3076.090 1810.310 3077.270 ;
        RECT 1810.730 3076.090 1811.910 3077.270 ;
        RECT 1809.130 3074.490 1810.310 3075.670 ;
        RECT 1810.730 3074.490 1811.910 3075.670 ;
        RECT 1809.130 2896.090 1810.310 2897.270 ;
        RECT 1810.730 2896.090 1811.910 2897.270 ;
        RECT 1809.130 2894.490 1810.310 2895.670 ;
        RECT 1810.730 2894.490 1811.910 2895.670 ;
        RECT 1809.130 2716.090 1810.310 2717.270 ;
        RECT 1810.730 2716.090 1811.910 2717.270 ;
        RECT 1809.130 2714.490 1810.310 2715.670 ;
        RECT 1810.730 2714.490 1811.910 2715.670 ;
        RECT 1809.130 2536.090 1810.310 2537.270 ;
        RECT 1810.730 2536.090 1811.910 2537.270 ;
        RECT 1809.130 2534.490 1810.310 2535.670 ;
        RECT 1810.730 2534.490 1811.910 2535.670 ;
        RECT 1809.130 2356.090 1810.310 2357.270 ;
        RECT 1810.730 2356.090 1811.910 2357.270 ;
        RECT 1809.130 2354.490 1810.310 2355.670 ;
        RECT 1810.730 2354.490 1811.910 2355.670 ;
        RECT 1809.130 2176.090 1810.310 2177.270 ;
        RECT 1810.730 2176.090 1811.910 2177.270 ;
        RECT 1809.130 2174.490 1810.310 2175.670 ;
        RECT 1810.730 2174.490 1811.910 2175.670 ;
        RECT 1809.130 1996.090 1810.310 1997.270 ;
        RECT 1810.730 1996.090 1811.910 1997.270 ;
        RECT 1809.130 1994.490 1810.310 1995.670 ;
        RECT 1810.730 1994.490 1811.910 1995.670 ;
        RECT 1809.130 1816.090 1810.310 1817.270 ;
        RECT 1810.730 1816.090 1811.910 1817.270 ;
        RECT 1809.130 1814.490 1810.310 1815.670 ;
        RECT 1810.730 1814.490 1811.910 1815.670 ;
        RECT 1809.130 1636.090 1810.310 1637.270 ;
        RECT 1810.730 1636.090 1811.910 1637.270 ;
        RECT 1809.130 1634.490 1810.310 1635.670 ;
        RECT 1810.730 1634.490 1811.910 1635.670 ;
        RECT 1809.130 1456.090 1810.310 1457.270 ;
        RECT 1810.730 1456.090 1811.910 1457.270 ;
        RECT 1809.130 1454.490 1810.310 1455.670 ;
        RECT 1810.730 1454.490 1811.910 1455.670 ;
        RECT 1809.130 1276.090 1810.310 1277.270 ;
        RECT 1810.730 1276.090 1811.910 1277.270 ;
        RECT 1809.130 1274.490 1810.310 1275.670 ;
        RECT 1810.730 1274.490 1811.910 1275.670 ;
        RECT 1809.130 1096.090 1810.310 1097.270 ;
        RECT 1810.730 1096.090 1811.910 1097.270 ;
        RECT 1809.130 1094.490 1810.310 1095.670 ;
        RECT 1810.730 1094.490 1811.910 1095.670 ;
        RECT 1809.130 916.090 1810.310 917.270 ;
        RECT 1810.730 916.090 1811.910 917.270 ;
        RECT 1809.130 914.490 1810.310 915.670 ;
        RECT 1810.730 914.490 1811.910 915.670 ;
        RECT 1809.130 736.090 1810.310 737.270 ;
        RECT 1810.730 736.090 1811.910 737.270 ;
        RECT 1809.130 734.490 1810.310 735.670 ;
        RECT 1810.730 734.490 1811.910 735.670 ;
        RECT 1809.130 556.090 1810.310 557.270 ;
        RECT 1810.730 556.090 1811.910 557.270 ;
        RECT 1809.130 554.490 1810.310 555.670 ;
        RECT 1810.730 554.490 1811.910 555.670 ;
        RECT 1809.130 376.090 1810.310 377.270 ;
        RECT 1810.730 376.090 1811.910 377.270 ;
        RECT 1809.130 374.490 1810.310 375.670 ;
        RECT 1810.730 374.490 1811.910 375.670 ;
        RECT 1809.130 196.090 1810.310 197.270 ;
        RECT 1810.730 196.090 1811.910 197.270 ;
        RECT 1809.130 194.490 1810.310 195.670 ;
        RECT 1810.730 194.490 1811.910 195.670 ;
        RECT 1809.130 16.090 1810.310 17.270 ;
        RECT 1810.730 16.090 1811.910 17.270 ;
        RECT 1809.130 14.490 1810.310 15.670 ;
        RECT 1810.730 14.490 1811.910 15.670 ;
        RECT 1809.130 -4.460 1810.310 -3.280 ;
        RECT 1810.730 -4.460 1811.910 -3.280 ;
        RECT 1809.130 -6.060 1810.310 -4.880 ;
        RECT 1810.730 -6.060 1811.910 -4.880 ;
        RECT 1989.130 3524.560 1990.310 3525.740 ;
        RECT 1990.730 3524.560 1991.910 3525.740 ;
        RECT 1989.130 3522.960 1990.310 3524.140 ;
        RECT 1990.730 3522.960 1991.910 3524.140 ;
        RECT 1989.130 3436.090 1990.310 3437.270 ;
        RECT 1990.730 3436.090 1991.910 3437.270 ;
        RECT 1989.130 3434.490 1990.310 3435.670 ;
        RECT 1990.730 3434.490 1991.910 3435.670 ;
        RECT 1989.130 3256.090 1990.310 3257.270 ;
        RECT 1990.730 3256.090 1991.910 3257.270 ;
        RECT 1989.130 3254.490 1990.310 3255.670 ;
        RECT 1990.730 3254.490 1991.910 3255.670 ;
        RECT 1989.130 3076.090 1990.310 3077.270 ;
        RECT 1990.730 3076.090 1991.910 3077.270 ;
        RECT 1989.130 3074.490 1990.310 3075.670 ;
        RECT 1990.730 3074.490 1991.910 3075.670 ;
        RECT 1989.130 2896.090 1990.310 2897.270 ;
        RECT 1990.730 2896.090 1991.910 2897.270 ;
        RECT 1989.130 2894.490 1990.310 2895.670 ;
        RECT 1990.730 2894.490 1991.910 2895.670 ;
        RECT 1989.130 2716.090 1990.310 2717.270 ;
        RECT 1990.730 2716.090 1991.910 2717.270 ;
        RECT 1989.130 2714.490 1990.310 2715.670 ;
        RECT 1990.730 2714.490 1991.910 2715.670 ;
        RECT 1989.130 2536.090 1990.310 2537.270 ;
        RECT 1990.730 2536.090 1991.910 2537.270 ;
        RECT 1989.130 2534.490 1990.310 2535.670 ;
        RECT 1990.730 2534.490 1991.910 2535.670 ;
        RECT 1989.130 2356.090 1990.310 2357.270 ;
        RECT 1990.730 2356.090 1991.910 2357.270 ;
        RECT 1989.130 2354.490 1990.310 2355.670 ;
        RECT 1990.730 2354.490 1991.910 2355.670 ;
        RECT 1989.130 2176.090 1990.310 2177.270 ;
        RECT 1990.730 2176.090 1991.910 2177.270 ;
        RECT 1989.130 2174.490 1990.310 2175.670 ;
        RECT 1990.730 2174.490 1991.910 2175.670 ;
        RECT 1989.130 1996.090 1990.310 1997.270 ;
        RECT 1990.730 1996.090 1991.910 1997.270 ;
        RECT 1989.130 1994.490 1990.310 1995.670 ;
        RECT 1990.730 1994.490 1991.910 1995.670 ;
        RECT 1989.130 1816.090 1990.310 1817.270 ;
        RECT 1990.730 1816.090 1991.910 1817.270 ;
        RECT 1989.130 1814.490 1990.310 1815.670 ;
        RECT 1990.730 1814.490 1991.910 1815.670 ;
        RECT 1989.130 1636.090 1990.310 1637.270 ;
        RECT 1990.730 1636.090 1991.910 1637.270 ;
        RECT 1989.130 1634.490 1990.310 1635.670 ;
        RECT 1990.730 1634.490 1991.910 1635.670 ;
        RECT 1989.130 1456.090 1990.310 1457.270 ;
        RECT 1990.730 1456.090 1991.910 1457.270 ;
        RECT 1989.130 1454.490 1990.310 1455.670 ;
        RECT 1990.730 1454.490 1991.910 1455.670 ;
        RECT 1989.130 1276.090 1990.310 1277.270 ;
        RECT 1990.730 1276.090 1991.910 1277.270 ;
        RECT 1989.130 1274.490 1990.310 1275.670 ;
        RECT 1990.730 1274.490 1991.910 1275.670 ;
        RECT 1989.130 1096.090 1990.310 1097.270 ;
        RECT 1990.730 1096.090 1991.910 1097.270 ;
        RECT 1989.130 1094.490 1990.310 1095.670 ;
        RECT 1990.730 1094.490 1991.910 1095.670 ;
        RECT 1989.130 916.090 1990.310 917.270 ;
        RECT 1990.730 916.090 1991.910 917.270 ;
        RECT 1989.130 914.490 1990.310 915.670 ;
        RECT 1990.730 914.490 1991.910 915.670 ;
        RECT 1989.130 736.090 1990.310 737.270 ;
        RECT 1990.730 736.090 1991.910 737.270 ;
        RECT 1989.130 734.490 1990.310 735.670 ;
        RECT 1990.730 734.490 1991.910 735.670 ;
        RECT 1989.130 556.090 1990.310 557.270 ;
        RECT 1990.730 556.090 1991.910 557.270 ;
        RECT 1989.130 554.490 1990.310 555.670 ;
        RECT 1990.730 554.490 1991.910 555.670 ;
        RECT 1989.130 376.090 1990.310 377.270 ;
        RECT 1990.730 376.090 1991.910 377.270 ;
        RECT 1989.130 374.490 1990.310 375.670 ;
        RECT 1990.730 374.490 1991.910 375.670 ;
        RECT 1989.130 196.090 1990.310 197.270 ;
        RECT 1990.730 196.090 1991.910 197.270 ;
        RECT 1989.130 194.490 1990.310 195.670 ;
        RECT 1990.730 194.490 1991.910 195.670 ;
        RECT 1989.130 16.090 1990.310 17.270 ;
        RECT 1990.730 16.090 1991.910 17.270 ;
        RECT 1989.130 14.490 1990.310 15.670 ;
        RECT 1990.730 14.490 1991.910 15.670 ;
        RECT 1989.130 -4.460 1990.310 -3.280 ;
        RECT 1990.730 -4.460 1991.910 -3.280 ;
        RECT 1989.130 -6.060 1990.310 -4.880 ;
        RECT 1990.730 -6.060 1991.910 -4.880 ;
        RECT 2169.130 3524.560 2170.310 3525.740 ;
        RECT 2170.730 3524.560 2171.910 3525.740 ;
        RECT 2169.130 3522.960 2170.310 3524.140 ;
        RECT 2170.730 3522.960 2171.910 3524.140 ;
        RECT 2169.130 3436.090 2170.310 3437.270 ;
        RECT 2170.730 3436.090 2171.910 3437.270 ;
        RECT 2169.130 3434.490 2170.310 3435.670 ;
        RECT 2170.730 3434.490 2171.910 3435.670 ;
        RECT 2169.130 3256.090 2170.310 3257.270 ;
        RECT 2170.730 3256.090 2171.910 3257.270 ;
        RECT 2169.130 3254.490 2170.310 3255.670 ;
        RECT 2170.730 3254.490 2171.910 3255.670 ;
        RECT 2169.130 3076.090 2170.310 3077.270 ;
        RECT 2170.730 3076.090 2171.910 3077.270 ;
        RECT 2169.130 3074.490 2170.310 3075.670 ;
        RECT 2170.730 3074.490 2171.910 3075.670 ;
        RECT 2169.130 2896.090 2170.310 2897.270 ;
        RECT 2170.730 2896.090 2171.910 2897.270 ;
        RECT 2169.130 2894.490 2170.310 2895.670 ;
        RECT 2170.730 2894.490 2171.910 2895.670 ;
        RECT 2169.130 2716.090 2170.310 2717.270 ;
        RECT 2170.730 2716.090 2171.910 2717.270 ;
        RECT 2169.130 2714.490 2170.310 2715.670 ;
        RECT 2170.730 2714.490 2171.910 2715.670 ;
        RECT 2169.130 2536.090 2170.310 2537.270 ;
        RECT 2170.730 2536.090 2171.910 2537.270 ;
        RECT 2169.130 2534.490 2170.310 2535.670 ;
        RECT 2170.730 2534.490 2171.910 2535.670 ;
        RECT 2169.130 2356.090 2170.310 2357.270 ;
        RECT 2170.730 2356.090 2171.910 2357.270 ;
        RECT 2169.130 2354.490 2170.310 2355.670 ;
        RECT 2170.730 2354.490 2171.910 2355.670 ;
        RECT 2169.130 2176.090 2170.310 2177.270 ;
        RECT 2170.730 2176.090 2171.910 2177.270 ;
        RECT 2169.130 2174.490 2170.310 2175.670 ;
        RECT 2170.730 2174.490 2171.910 2175.670 ;
        RECT 2169.130 1996.090 2170.310 1997.270 ;
        RECT 2170.730 1996.090 2171.910 1997.270 ;
        RECT 2169.130 1994.490 2170.310 1995.670 ;
        RECT 2170.730 1994.490 2171.910 1995.670 ;
        RECT 2169.130 1816.090 2170.310 1817.270 ;
        RECT 2170.730 1816.090 2171.910 1817.270 ;
        RECT 2169.130 1814.490 2170.310 1815.670 ;
        RECT 2170.730 1814.490 2171.910 1815.670 ;
        RECT 2169.130 1636.090 2170.310 1637.270 ;
        RECT 2170.730 1636.090 2171.910 1637.270 ;
        RECT 2169.130 1634.490 2170.310 1635.670 ;
        RECT 2170.730 1634.490 2171.910 1635.670 ;
        RECT 2169.130 1456.090 2170.310 1457.270 ;
        RECT 2170.730 1456.090 2171.910 1457.270 ;
        RECT 2169.130 1454.490 2170.310 1455.670 ;
        RECT 2170.730 1454.490 2171.910 1455.670 ;
        RECT 2169.130 1276.090 2170.310 1277.270 ;
        RECT 2170.730 1276.090 2171.910 1277.270 ;
        RECT 2169.130 1274.490 2170.310 1275.670 ;
        RECT 2170.730 1274.490 2171.910 1275.670 ;
        RECT 2169.130 1096.090 2170.310 1097.270 ;
        RECT 2170.730 1096.090 2171.910 1097.270 ;
        RECT 2169.130 1094.490 2170.310 1095.670 ;
        RECT 2170.730 1094.490 2171.910 1095.670 ;
        RECT 2169.130 916.090 2170.310 917.270 ;
        RECT 2170.730 916.090 2171.910 917.270 ;
        RECT 2169.130 914.490 2170.310 915.670 ;
        RECT 2170.730 914.490 2171.910 915.670 ;
        RECT 2169.130 736.090 2170.310 737.270 ;
        RECT 2170.730 736.090 2171.910 737.270 ;
        RECT 2169.130 734.490 2170.310 735.670 ;
        RECT 2170.730 734.490 2171.910 735.670 ;
        RECT 2169.130 556.090 2170.310 557.270 ;
        RECT 2170.730 556.090 2171.910 557.270 ;
        RECT 2169.130 554.490 2170.310 555.670 ;
        RECT 2170.730 554.490 2171.910 555.670 ;
        RECT 2169.130 376.090 2170.310 377.270 ;
        RECT 2170.730 376.090 2171.910 377.270 ;
        RECT 2169.130 374.490 2170.310 375.670 ;
        RECT 2170.730 374.490 2171.910 375.670 ;
        RECT 2169.130 196.090 2170.310 197.270 ;
        RECT 2170.730 196.090 2171.910 197.270 ;
        RECT 2169.130 194.490 2170.310 195.670 ;
        RECT 2170.730 194.490 2171.910 195.670 ;
        RECT 2169.130 16.090 2170.310 17.270 ;
        RECT 2170.730 16.090 2171.910 17.270 ;
        RECT 2169.130 14.490 2170.310 15.670 ;
        RECT 2170.730 14.490 2171.910 15.670 ;
        RECT 2169.130 -4.460 2170.310 -3.280 ;
        RECT 2170.730 -4.460 2171.910 -3.280 ;
        RECT 2169.130 -6.060 2170.310 -4.880 ;
        RECT 2170.730 -6.060 2171.910 -4.880 ;
        RECT 2349.130 3524.560 2350.310 3525.740 ;
        RECT 2350.730 3524.560 2351.910 3525.740 ;
        RECT 2349.130 3522.960 2350.310 3524.140 ;
        RECT 2350.730 3522.960 2351.910 3524.140 ;
        RECT 2349.130 3436.090 2350.310 3437.270 ;
        RECT 2350.730 3436.090 2351.910 3437.270 ;
        RECT 2349.130 3434.490 2350.310 3435.670 ;
        RECT 2350.730 3434.490 2351.910 3435.670 ;
        RECT 2349.130 3256.090 2350.310 3257.270 ;
        RECT 2350.730 3256.090 2351.910 3257.270 ;
        RECT 2349.130 3254.490 2350.310 3255.670 ;
        RECT 2350.730 3254.490 2351.910 3255.670 ;
        RECT 2349.130 3076.090 2350.310 3077.270 ;
        RECT 2350.730 3076.090 2351.910 3077.270 ;
        RECT 2349.130 3074.490 2350.310 3075.670 ;
        RECT 2350.730 3074.490 2351.910 3075.670 ;
        RECT 2349.130 2896.090 2350.310 2897.270 ;
        RECT 2350.730 2896.090 2351.910 2897.270 ;
        RECT 2349.130 2894.490 2350.310 2895.670 ;
        RECT 2350.730 2894.490 2351.910 2895.670 ;
        RECT 2349.130 2716.090 2350.310 2717.270 ;
        RECT 2350.730 2716.090 2351.910 2717.270 ;
        RECT 2349.130 2714.490 2350.310 2715.670 ;
        RECT 2350.730 2714.490 2351.910 2715.670 ;
        RECT 2349.130 2536.090 2350.310 2537.270 ;
        RECT 2350.730 2536.090 2351.910 2537.270 ;
        RECT 2349.130 2534.490 2350.310 2535.670 ;
        RECT 2350.730 2534.490 2351.910 2535.670 ;
        RECT 2349.130 2356.090 2350.310 2357.270 ;
        RECT 2350.730 2356.090 2351.910 2357.270 ;
        RECT 2349.130 2354.490 2350.310 2355.670 ;
        RECT 2350.730 2354.490 2351.910 2355.670 ;
        RECT 2349.130 2176.090 2350.310 2177.270 ;
        RECT 2350.730 2176.090 2351.910 2177.270 ;
        RECT 2349.130 2174.490 2350.310 2175.670 ;
        RECT 2350.730 2174.490 2351.910 2175.670 ;
        RECT 2349.130 1996.090 2350.310 1997.270 ;
        RECT 2350.730 1996.090 2351.910 1997.270 ;
        RECT 2349.130 1994.490 2350.310 1995.670 ;
        RECT 2350.730 1994.490 2351.910 1995.670 ;
        RECT 2349.130 1816.090 2350.310 1817.270 ;
        RECT 2350.730 1816.090 2351.910 1817.270 ;
        RECT 2349.130 1814.490 2350.310 1815.670 ;
        RECT 2350.730 1814.490 2351.910 1815.670 ;
        RECT 2349.130 1636.090 2350.310 1637.270 ;
        RECT 2350.730 1636.090 2351.910 1637.270 ;
        RECT 2349.130 1634.490 2350.310 1635.670 ;
        RECT 2350.730 1634.490 2351.910 1635.670 ;
        RECT 2349.130 1456.090 2350.310 1457.270 ;
        RECT 2350.730 1456.090 2351.910 1457.270 ;
        RECT 2349.130 1454.490 2350.310 1455.670 ;
        RECT 2350.730 1454.490 2351.910 1455.670 ;
        RECT 2349.130 1276.090 2350.310 1277.270 ;
        RECT 2350.730 1276.090 2351.910 1277.270 ;
        RECT 2349.130 1274.490 2350.310 1275.670 ;
        RECT 2350.730 1274.490 2351.910 1275.670 ;
        RECT 2349.130 1096.090 2350.310 1097.270 ;
        RECT 2350.730 1096.090 2351.910 1097.270 ;
        RECT 2349.130 1094.490 2350.310 1095.670 ;
        RECT 2350.730 1094.490 2351.910 1095.670 ;
        RECT 2349.130 916.090 2350.310 917.270 ;
        RECT 2350.730 916.090 2351.910 917.270 ;
        RECT 2349.130 914.490 2350.310 915.670 ;
        RECT 2350.730 914.490 2351.910 915.670 ;
        RECT 2349.130 736.090 2350.310 737.270 ;
        RECT 2350.730 736.090 2351.910 737.270 ;
        RECT 2349.130 734.490 2350.310 735.670 ;
        RECT 2350.730 734.490 2351.910 735.670 ;
        RECT 2349.130 556.090 2350.310 557.270 ;
        RECT 2350.730 556.090 2351.910 557.270 ;
        RECT 2349.130 554.490 2350.310 555.670 ;
        RECT 2350.730 554.490 2351.910 555.670 ;
        RECT 2349.130 376.090 2350.310 377.270 ;
        RECT 2350.730 376.090 2351.910 377.270 ;
        RECT 2349.130 374.490 2350.310 375.670 ;
        RECT 2350.730 374.490 2351.910 375.670 ;
        RECT 2349.130 196.090 2350.310 197.270 ;
        RECT 2350.730 196.090 2351.910 197.270 ;
        RECT 2349.130 194.490 2350.310 195.670 ;
        RECT 2350.730 194.490 2351.910 195.670 ;
        RECT 2349.130 16.090 2350.310 17.270 ;
        RECT 2350.730 16.090 2351.910 17.270 ;
        RECT 2349.130 14.490 2350.310 15.670 ;
        RECT 2350.730 14.490 2351.910 15.670 ;
        RECT 2349.130 -4.460 2350.310 -3.280 ;
        RECT 2350.730 -4.460 2351.910 -3.280 ;
        RECT 2349.130 -6.060 2350.310 -4.880 ;
        RECT 2350.730 -6.060 2351.910 -4.880 ;
        RECT 2529.130 3524.560 2530.310 3525.740 ;
        RECT 2530.730 3524.560 2531.910 3525.740 ;
        RECT 2529.130 3522.960 2530.310 3524.140 ;
        RECT 2530.730 3522.960 2531.910 3524.140 ;
        RECT 2529.130 3436.090 2530.310 3437.270 ;
        RECT 2530.730 3436.090 2531.910 3437.270 ;
        RECT 2529.130 3434.490 2530.310 3435.670 ;
        RECT 2530.730 3434.490 2531.910 3435.670 ;
        RECT 2529.130 3256.090 2530.310 3257.270 ;
        RECT 2530.730 3256.090 2531.910 3257.270 ;
        RECT 2529.130 3254.490 2530.310 3255.670 ;
        RECT 2530.730 3254.490 2531.910 3255.670 ;
        RECT 2529.130 3076.090 2530.310 3077.270 ;
        RECT 2530.730 3076.090 2531.910 3077.270 ;
        RECT 2529.130 3074.490 2530.310 3075.670 ;
        RECT 2530.730 3074.490 2531.910 3075.670 ;
        RECT 2529.130 2896.090 2530.310 2897.270 ;
        RECT 2530.730 2896.090 2531.910 2897.270 ;
        RECT 2529.130 2894.490 2530.310 2895.670 ;
        RECT 2530.730 2894.490 2531.910 2895.670 ;
        RECT 2529.130 2716.090 2530.310 2717.270 ;
        RECT 2530.730 2716.090 2531.910 2717.270 ;
        RECT 2529.130 2714.490 2530.310 2715.670 ;
        RECT 2530.730 2714.490 2531.910 2715.670 ;
        RECT 2529.130 2536.090 2530.310 2537.270 ;
        RECT 2530.730 2536.090 2531.910 2537.270 ;
        RECT 2529.130 2534.490 2530.310 2535.670 ;
        RECT 2530.730 2534.490 2531.910 2535.670 ;
        RECT 2529.130 2356.090 2530.310 2357.270 ;
        RECT 2530.730 2356.090 2531.910 2357.270 ;
        RECT 2529.130 2354.490 2530.310 2355.670 ;
        RECT 2530.730 2354.490 2531.910 2355.670 ;
        RECT 2529.130 2176.090 2530.310 2177.270 ;
        RECT 2530.730 2176.090 2531.910 2177.270 ;
        RECT 2529.130 2174.490 2530.310 2175.670 ;
        RECT 2530.730 2174.490 2531.910 2175.670 ;
        RECT 2529.130 1996.090 2530.310 1997.270 ;
        RECT 2530.730 1996.090 2531.910 1997.270 ;
        RECT 2529.130 1994.490 2530.310 1995.670 ;
        RECT 2530.730 1994.490 2531.910 1995.670 ;
        RECT 2529.130 1816.090 2530.310 1817.270 ;
        RECT 2530.730 1816.090 2531.910 1817.270 ;
        RECT 2529.130 1814.490 2530.310 1815.670 ;
        RECT 2530.730 1814.490 2531.910 1815.670 ;
        RECT 2529.130 1636.090 2530.310 1637.270 ;
        RECT 2530.730 1636.090 2531.910 1637.270 ;
        RECT 2529.130 1634.490 2530.310 1635.670 ;
        RECT 2530.730 1634.490 2531.910 1635.670 ;
        RECT 2529.130 1456.090 2530.310 1457.270 ;
        RECT 2530.730 1456.090 2531.910 1457.270 ;
        RECT 2529.130 1454.490 2530.310 1455.670 ;
        RECT 2530.730 1454.490 2531.910 1455.670 ;
        RECT 2529.130 1276.090 2530.310 1277.270 ;
        RECT 2530.730 1276.090 2531.910 1277.270 ;
        RECT 2529.130 1274.490 2530.310 1275.670 ;
        RECT 2530.730 1274.490 2531.910 1275.670 ;
        RECT 2529.130 1096.090 2530.310 1097.270 ;
        RECT 2530.730 1096.090 2531.910 1097.270 ;
        RECT 2529.130 1094.490 2530.310 1095.670 ;
        RECT 2530.730 1094.490 2531.910 1095.670 ;
        RECT 2529.130 916.090 2530.310 917.270 ;
        RECT 2530.730 916.090 2531.910 917.270 ;
        RECT 2529.130 914.490 2530.310 915.670 ;
        RECT 2530.730 914.490 2531.910 915.670 ;
        RECT 2529.130 736.090 2530.310 737.270 ;
        RECT 2530.730 736.090 2531.910 737.270 ;
        RECT 2529.130 734.490 2530.310 735.670 ;
        RECT 2530.730 734.490 2531.910 735.670 ;
        RECT 2529.130 556.090 2530.310 557.270 ;
        RECT 2530.730 556.090 2531.910 557.270 ;
        RECT 2529.130 554.490 2530.310 555.670 ;
        RECT 2530.730 554.490 2531.910 555.670 ;
        RECT 2529.130 376.090 2530.310 377.270 ;
        RECT 2530.730 376.090 2531.910 377.270 ;
        RECT 2529.130 374.490 2530.310 375.670 ;
        RECT 2530.730 374.490 2531.910 375.670 ;
        RECT 2529.130 196.090 2530.310 197.270 ;
        RECT 2530.730 196.090 2531.910 197.270 ;
        RECT 2529.130 194.490 2530.310 195.670 ;
        RECT 2530.730 194.490 2531.910 195.670 ;
        RECT 2529.130 16.090 2530.310 17.270 ;
        RECT 2530.730 16.090 2531.910 17.270 ;
        RECT 2529.130 14.490 2530.310 15.670 ;
        RECT 2530.730 14.490 2531.910 15.670 ;
        RECT 2529.130 -4.460 2530.310 -3.280 ;
        RECT 2530.730 -4.460 2531.910 -3.280 ;
        RECT 2529.130 -6.060 2530.310 -4.880 ;
        RECT 2530.730 -6.060 2531.910 -4.880 ;
        RECT 2709.130 3524.560 2710.310 3525.740 ;
        RECT 2710.730 3524.560 2711.910 3525.740 ;
        RECT 2709.130 3522.960 2710.310 3524.140 ;
        RECT 2710.730 3522.960 2711.910 3524.140 ;
        RECT 2709.130 3436.090 2710.310 3437.270 ;
        RECT 2710.730 3436.090 2711.910 3437.270 ;
        RECT 2709.130 3434.490 2710.310 3435.670 ;
        RECT 2710.730 3434.490 2711.910 3435.670 ;
        RECT 2709.130 3256.090 2710.310 3257.270 ;
        RECT 2710.730 3256.090 2711.910 3257.270 ;
        RECT 2709.130 3254.490 2710.310 3255.670 ;
        RECT 2710.730 3254.490 2711.910 3255.670 ;
        RECT 2709.130 3076.090 2710.310 3077.270 ;
        RECT 2710.730 3076.090 2711.910 3077.270 ;
        RECT 2709.130 3074.490 2710.310 3075.670 ;
        RECT 2710.730 3074.490 2711.910 3075.670 ;
        RECT 2709.130 2896.090 2710.310 2897.270 ;
        RECT 2710.730 2896.090 2711.910 2897.270 ;
        RECT 2709.130 2894.490 2710.310 2895.670 ;
        RECT 2710.730 2894.490 2711.910 2895.670 ;
        RECT 2709.130 2716.090 2710.310 2717.270 ;
        RECT 2710.730 2716.090 2711.910 2717.270 ;
        RECT 2709.130 2714.490 2710.310 2715.670 ;
        RECT 2710.730 2714.490 2711.910 2715.670 ;
        RECT 2709.130 2536.090 2710.310 2537.270 ;
        RECT 2710.730 2536.090 2711.910 2537.270 ;
        RECT 2709.130 2534.490 2710.310 2535.670 ;
        RECT 2710.730 2534.490 2711.910 2535.670 ;
        RECT 2709.130 2356.090 2710.310 2357.270 ;
        RECT 2710.730 2356.090 2711.910 2357.270 ;
        RECT 2709.130 2354.490 2710.310 2355.670 ;
        RECT 2710.730 2354.490 2711.910 2355.670 ;
        RECT 2709.130 2176.090 2710.310 2177.270 ;
        RECT 2710.730 2176.090 2711.910 2177.270 ;
        RECT 2709.130 2174.490 2710.310 2175.670 ;
        RECT 2710.730 2174.490 2711.910 2175.670 ;
        RECT 2709.130 1996.090 2710.310 1997.270 ;
        RECT 2710.730 1996.090 2711.910 1997.270 ;
        RECT 2709.130 1994.490 2710.310 1995.670 ;
        RECT 2710.730 1994.490 2711.910 1995.670 ;
        RECT 2709.130 1816.090 2710.310 1817.270 ;
        RECT 2710.730 1816.090 2711.910 1817.270 ;
        RECT 2709.130 1814.490 2710.310 1815.670 ;
        RECT 2710.730 1814.490 2711.910 1815.670 ;
        RECT 2709.130 1636.090 2710.310 1637.270 ;
        RECT 2710.730 1636.090 2711.910 1637.270 ;
        RECT 2709.130 1634.490 2710.310 1635.670 ;
        RECT 2710.730 1634.490 2711.910 1635.670 ;
        RECT 2709.130 1456.090 2710.310 1457.270 ;
        RECT 2710.730 1456.090 2711.910 1457.270 ;
        RECT 2709.130 1454.490 2710.310 1455.670 ;
        RECT 2710.730 1454.490 2711.910 1455.670 ;
        RECT 2709.130 1276.090 2710.310 1277.270 ;
        RECT 2710.730 1276.090 2711.910 1277.270 ;
        RECT 2709.130 1274.490 2710.310 1275.670 ;
        RECT 2710.730 1274.490 2711.910 1275.670 ;
        RECT 2709.130 1096.090 2710.310 1097.270 ;
        RECT 2710.730 1096.090 2711.910 1097.270 ;
        RECT 2709.130 1094.490 2710.310 1095.670 ;
        RECT 2710.730 1094.490 2711.910 1095.670 ;
        RECT 2709.130 916.090 2710.310 917.270 ;
        RECT 2710.730 916.090 2711.910 917.270 ;
        RECT 2709.130 914.490 2710.310 915.670 ;
        RECT 2710.730 914.490 2711.910 915.670 ;
        RECT 2709.130 736.090 2710.310 737.270 ;
        RECT 2710.730 736.090 2711.910 737.270 ;
        RECT 2709.130 734.490 2710.310 735.670 ;
        RECT 2710.730 734.490 2711.910 735.670 ;
        RECT 2709.130 556.090 2710.310 557.270 ;
        RECT 2710.730 556.090 2711.910 557.270 ;
        RECT 2709.130 554.490 2710.310 555.670 ;
        RECT 2710.730 554.490 2711.910 555.670 ;
        RECT 2709.130 376.090 2710.310 377.270 ;
        RECT 2710.730 376.090 2711.910 377.270 ;
        RECT 2709.130 374.490 2710.310 375.670 ;
        RECT 2710.730 374.490 2711.910 375.670 ;
        RECT 2709.130 196.090 2710.310 197.270 ;
        RECT 2710.730 196.090 2711.910 197.270 ;
        RECT 2709.130 194.490 2710.310 195.670 ;
        RECT 2710.730 194.490 2711.910 195.670 ;
        RECT 2709.130 16.090 2710.310 17.270 ;
        RECT 2710.730 16.090 2711.910 17.270 ;
        RECT 2709.130 14.490 2710.310 15.670 ;
        RECT 2710.730 14.490 2711.910 15.670 ;
        RECT 2709.130 -4.460 2710.310 -3.280 ;
        RECT 2710.730 -4.460 2711.910 -3.280 ;
        RECT 2709.130 -6.060 2710.310 -4.880 ;
        RECT 2710.730 -6.060 2711.910 -4.880 ;
        RECT 2889.130 3524.560 2890.310 3525.740 ;
        RECT 2890.730 3524.560 2891.910 3525.740 ;
        RECT 2889.130 3522.960 2890.310 3524.140 ;
        RECT 2890.730 3522.960 2891.910 3524.140 ;
        RECT 2889.130 3436.090 2890.310 3437.270 ;
        RECT 2890.730 3436.090 2891.910 3437.270 ;
        RECT 2889.130 3434.490 2890.310 3435.670 ;
        RECT 2890.730 3434.490 2891.910 3435.670 ;
        RECT 2889.130 3256.090 2890.310 3257.270 ;
        RECT 2890.730 3256.090 2891.910 3257.270 ;
        RECT 2889.130 3254.490 2890.310 3255.670 ;
        RECT 2890.730 3254.490 2891.910 3255.670 ;
        RECT 2889.130 3076.090 2890.310 3077.270 ;
        RECT 2890.730 3076.090 2891.910 3077.270 ;
        RECT 2889.130 3074.490 2890.310 3075.670 ;
        RECT 2890.730 3074.490 2891.910 3075.670 ;
        RECT 2889.130 2896.090 2890.310 2897.270 ;
        RECT 2890.730 2896.090 2891.910 2897.270 ;
        RECT 2889.130 2894.490 2890.310 2895.670 ;
        RECT 2890.730 2894.490 2891.910 2895.670 ;
        RECT 2889.130 2716.090 2890.310 2717.270 ;
        RECT 2890.730 2716.090 2891.910 2717.270 ;
        RECT 2889.130 2714.490 2890.310 2715.670 ;
        RECT 2890.730 2714.490 2891.910 2715.670 ;
        RECT 2889.130 2536.090 2890.310 2537.270 ;
        RECT 2890.730 2536.090 2891.910 2537.270 ;
        RECT 2889.130 2534.490 2890.310 2535.670 ;
        RECT 2890.730 2534.490 2891.910 2535.670 ;
        RECT 2889.130 2356.090 2890.310 2357.270 ;
        RECT 2890.730 2356.090 2891.910 2357.270 ;
        RECT 2889.130 2354.490 2890.310 2355.670 ;
        RECT 2890.730 2354.490 2891.910 2355.670 ;
        RECT 2889.130 2176.090 2890.310 2177.270 ;
        RECT 2890.730 2176.090 2891.910 2177.270 ;
        RECT 2889.130 2174.490 2890.310 2175.670 ;
        RECT 2890.730 2174.490 2891.910 2175.670 ;
        RECT 2889.130 1996.090 2890.310 1997.270 ;
        RECT 2890.730 1996.090 2891.910 1997.270 ;
        RECT 2889.130 1994.490 2890.310 1995.670 ;
        RECT 2890.730 1994.490 2891.910 1995.670 ;
        RECT 2889.130 1816.090 2890.310 1817.270 ;
        RECT 2890.730 1816.090 2891.910 1817.270 ;
        RECT 2889.130 1814.490 2890.310 1815.670 ;
        RECT 2890.730 1814.490 2891.910 1815.670 ;
        RECT 2889.130 1636.090 2890.310 1637.270 ;
        RECT 2890.730 1636.090 2891.910 1637.270 ;
        RECT 2889.130 1634.490 2890.310 1635.670 ;
        RECT 2890.730 1634.490 2891.910 1635.670 ;
        RECT 2889.130 1456.090 2890.310 1457.270 ;
        RECT 2890.730 1456.090 2891.910 1457.270 ;
        RECT 2889.130 1454.490 2890.310 1455.670 ;
        RECT 2890.730 1454.490 2891.910 1455.670 ;
        RECT 2889.130 1276.090 2890.310 1277.270 ;
        RECT 2890.730 1276.090 2891.910 1277.270 ;
        RECT 2889.130 1274.490 2890.310 1275.670 ;
        RECT 2890.730 1274.490 2891.910 1275.670 ;
        RECT 2889.130 1096.090 2890.310 1097.270 ;
        RECT 2890.730 1096.090 2891.910 1097.270 ;
        RECT 2889.130 1094.490 2890.310 1095.670 ;
        RECT 2890.730 1094.490 2891.910 1095.670 ;
        RECT 2889.130 916.090 2890.310 917.270 ;
        RECT 2890.730 916.090 2891.910 917.270 ;
        RECT 2889.130 914.490 2890.310 915.670 ;
        RECT 2890.730 914.490 2891.910 915.670 ;
        RECT 2889.130 736.090 2890.310 737.270 ;
        RECT 2890.730 736.090 2891.910 737.270 ;
        RECT 2889.130 734.490 2890.310 735.670 ;
        RECT 2890.730 734.490 2891.910 735.670 ;
        RECT 2889.130 556.090 2890.310 557.270 ;
        RECT 2890.730 556.090 2891.910 557.270 ;
        RECT 2889.130 554.490 2890.310 555.670 ;
        RECT 2890.730 554.490 2891.910 555.670 ;
        RECT 2889.130 376.090 2890.310 377.270 ;
        RECT 2890.730 376.090 2891.910 377.270 ;
        RECT 2889.130 374.490 2890.310 375.670 ;
        RECT 2890.730 374.490 2891.910 375.670 ;
        RECT 2889.130 196.090 2890.310 197.270 ;
        RECT 2890.730 196.090 2891.910 197.270 ;
        RECT 2889.130 194.490 2890.310 195.670 ;
        RECT 2890.730 194.490 2891.910 195.670 ;
        RECT 2889.130 16.090 2890.310 17.270 ;
        RECT 2890.730 16.090 2891.910 17.270 ;
        RECT 2889.130 14.490 2890.310 15.670 ;
        RECT 2890.730 14.490 2891.910 15.670 ;
        RECT 2889.130 -4.460 2890.310 -3.280 ;
        RECT 2890.730 -4.460 2891.910 -3.280 ;
        RECT 2889.130 -6.060 2890.310 -4.880 ;
        RECT 2890.730 -6.060 2891.910 -4.880 ;
        RECT 2928.260 3524.560 2929.440 3525.740 ;
        RECT 2929.860 3524.560 2931.040 3525.740 ;
        RECT 2928.260 3522.960 2929.440 3524.140 ;
        RECT 2929.860 3522.960 2931.040 3524.140 ;
        RECT 2928.260 3436.090 2929.440 3437.270 ;
        RECT 2929.860 3436.090 2931.040 3437.270 ;
        RECT 2928.260 3434.490 2929.440 3435.670 ;
        RECT 2929.860 3434.490 2931.040 3435.670 ;
        RECT 2928.260 3256.090 2929.440 3257.270 ;
        RECT 2929.860 3256.090 2931.040 3257.270 ;
        RECT 2928.260 3254.490 2929.440 3255.670 ;
        RECT 2929.860 3254.490 2931.040 3255.670 ;
        RECT 2928.260 3076.090 2929.440 3077.270 ;
        RECT 2929.860 3076.090 2931.040 3077.270 ;
        RECT 2928.260 3074.490 2929.440 3075.670 ;
        RECT 2929.860 3074.490 2931.040 3075.670 ;
        RECT 2928.260 2896.090 2929.440 2897.270 ;
        RECT 2929.860 2896.090 2931.040 2897.270 ;
        RECT 2928.260 2894.490 2929.440 2895.670 ;
        RECT 2929.860 2894.490 2931.040 2895.670 ;
        RECT 2928.260 2716.090 2929.440 2717.270 ;
        RECT 2929.860 2716.090 2931.040 2717.270 ;
        RECT 2928.260 2714.490 2929.440 2715.670 ;
        RECT 2929.860 2714.490 2931.040 2715.670 ;
        RECT 2928.260 2536.090 2929.440 2537.270 ;
        RECT 2929.860 2536.090 2931.040 2537.270 ;
        RECT 2928.260 2534.490 2929.440 2535.670 ;
        RECT 2929.860 2534.490 2931.040 2535.670 ;
        RECT 2928.260 2356.090 2929.440 2357.270 ;
        RECT 2929.860 2356.090 2931.040 2357.270 ;
        RECT 2928.260 2354.490 2929.440 2355.670 ;
        RECT 2929.860 2354.490 2931.040 2355.670 ;
        RECT 2928.260 2176.090 2929.440 2177.270 ;
        RECT 2929.860 2176.090 2931.040 2177.270 ;
        RECT 2928.260 2174.490 2929.440 2175.670 ;
        RECT 2929.860 2174.490 2931.040 2175.670 ;
        RECT 2928.260 1996.090 2929.440 1997.270 ;
        RECT 2929.860 1996.090 2931.040 1997.270 ;
        RECT 2928.260 1994.490 2929.440 1995.670 ;
        RECT 2929.860 1994.490 2931.040 1995.670 ;
        RECT 2928.260 1816.090 2929.440 1817.270 ;
        RECT 2929.860 1816.090 2931.040 1817.270 ;
        RECT 2928.260 1814.490 2929.440 1815.670 ;
        RECT 2929.860 1814.490 2931.040 1815.670 ;
        RECT 2928.260 1636.090 2929.440 1637.270 ;
        RECT 2929.860 1636.090 2931.040 1637.270 ;
        RECT 2928.260 1634.490 2929.440 1635.670 ;
        RECT 2929.860 1634.490 2931.040 1635.670 ;
        RECT 2928.260 1456.090 2929.440 1457.270 ;
        RECT 2929.860 1456.090 2931.040 1457.270 ;
        RECT 2928.260 1454.490 2929.440 1455.670 ;
        RECT 2929.860 1454.490 2931.040 1455.670 ;
        RECT 2928.260 1276.090 2929.440 1277.270 ;
        RECT 2929.860 1276.090 2931.040 1277.270 ;
        RECT 2928.260 1274.490 2929.440 1275.670 ;
        RECT 2929.860 1274.490 2931.040 1275.670 ;
        RECT 2928.260 1096.090 2929.440 1097.270 ;
        RECT 2929.860 1096.090 2931.040 1097.270 ;
        RECT 2928.260 1094.490 2929.440 1095.670 ;
        RECT 2929.860 1094.490 2931.040 1095.670 ;
        RECT 2928.260 916.090 2929.440 917.270 ;
        RECT 2929.860 916.090 2931.040 917.270 ;
        RECT 2928.260 914.490 2929.440 915.670 ;
        RECT 2929.860 914.490 2931.040 915.670 ;
        RECT 2928.260 736.090 2929.440 737.270 ;
        RECT 2929.860 736.090 2931.040 737.270 ;
        RECT 2928.260 734.490 2929.440 735.670 ;
        RECT 2929.860 734.490 2931.040 735.670 ;
        RECT 2928.260 556.090 2929.440 557.270 ;
        RECT 2929.860 556.090 2931.040 557.270 ;
        RECT 2928.260 554.490 2929.440 555.670 ;
        RECT 2929.860 554.490 2931.040 555.670 ;
        RECT 2928.260 376.090 2929.440 377.270 ;
        RECT 2929.860 376.090 2931.040 377.270 ;
        RECT 2928.260 374.490 2929.440 375.670 ;
        RECT 2929.860 374.490 2931.040 375.670 ;
        RECT 2928.260 196.090 2929.440 197.270 ;
        RECT 2929.860 196.090 2931.040 197.270 ;
        RECT 2928.260 194.490 2929.440 195.670 ;
        RECT 2929.860 194.490 2931.040 195.670 ;
        RECT 2928.260 16.090 2929.440 17.270 ;
        RECT 2929.860 16.090 2931.040 17.270 ;
        RECT 2928.260 14.490 2929.440 15.670 ;
        RECT 2929.860 14.490 2931.040 15.670 ;
        RECT 2928.260 -4.460 2929.440 -3.280 ;
        RECT 2929.860 -4.460 2931.040 -3.280 ;
        RECT 2928.260 -6.060 2929.440 -4.880 ;
        RECT 2929.860 -6.060 2931.040 -4.880 ;
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
        RECT -45.180 3434.330 2964.800 3437.430 ;
        RECT -45.180 3254.330 2964.800 3257.430 ;
        RECT -45.180 3074.330 2964.800 3077.430 ;
        RECT -45.180 2894.330 2964.800 2897.430 ;
        RECT -45.180 2714.330 2964.800 2717.430 ;
        RECT -45.180 2534.330 2964.800 2537.430 ;
        RECT -45.180 2354.330 2964.800 2357.430 ;
        RECT -45.180 2174.330 2964.800 2177.430 ;
        RECT -45.180 1994.330 2964.800 1997.430 ;
        RECT -45.180 1814.330 2964.800 1817.430 ;
        RECT -45.180 1634.330 2964.800 1637.430 ;
        RECT -45.180 1454.330 2964.800 1457.430 ;
        RECT -45.180 1274.330 2964.800 1277.430 ;
        RECT -45.180 1094.330 2964.800 1097.430 ;
        RECT -45.180 914.330 2964.800 917.430 ;
        RECT -45.180 734.330 2964.800 737.430 ;
        RECT -45.180 554.330 2964.800 557.430 ;
        RECT -45.180 374.330 2964.800 377.430 ;
        RECT -45.180 194.330 2964.800 197.430 ;
        RECT -45.180 14.330 2964.800 17.430 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -21.180 -15.820 -18.080 3535.500 ;
        RECT 53.970 -39.820 57.070 3559.500 ;
        RECT 233.970 -39.820 237.070 3559.500 ;
        RECT 413.970 760.000 417.070 3559.500 ;
        RECT 593.970 760.000 597.070 3559.500 ;
        RECT 413.970 -39.820 417.070 490.000 ;
        RECT 593.970 -39.820 597.070 490.000 ;
        RECT 773.970 -39.820 777.070 3559.500 ;
        RECT 953.970 -39.820 957.070 3559.500 ;
        RECT 1133.970 -39.820 1137.070 3559.500 ;
        RECT 1313.970 -39.820 1317.070 3559.500 ;
        RECT 1493.970 -39.820 1497.070 3559.500 ;
        RECT 1673.970 -39.820 1677.070 3559.500 ;
        RECT 1853.970 -39.820 1857.070 3559.500 ;
        RECT 2033.970 -39.820 2037.070 3559.500 ;
        RECT 2213.970 -39.820 2217.070 3559.500 ;
        RECT 2393.970 -39.820 2397.070 3559.500 ;
        RECT 2573.970 -39.820 2577.070 3559.500 ;
        RECT 2753.970 -39.820 2757.070 3559.500 ;
        RECT 2937.700 -15.820 2940.800 3535.500 ;
      LAYER via4 ;
        RECT -21.020 3534.160 -19.840 3535.340 ;
        RECT -19.420 3534.160 -18.240 3535.340 ;
        RECT -21.020 3532.560 -19.840 3533.740 ;
        RECT -19.420 3532.560 -18.240 3533.740 ;
        RECT -21.020 3481.090 -19.840 3482.270 ;
        RECT -19.420 3481.090 -18.240 3482.270 ;
        RECT -21.020 3479.490 -19.840 3480.670 ;
        RECT -19.420 3479.490 -18.240 3480.670 ;
        RECT -21.020 3301.090 -19.840 3302.270 ;
        RECT -19.420 3301.090 -18.240 3302.270 ;
        RECT -21.020 3299.490 -19.840 3300.670 ;
        RECT -19.420 3299.490 -18.240 3300.670 ;
        RECT -21.020 3121.090 -19.840 3122.270 ;
        RECT -19.420 3121.090 -18.240 3122.270 ;
        RECT -21.020 3119.490 -19.840 3120.670 ;
        RECT -19.420 3119.490 -18.240 3120.670 ;
        RECT -21.020 2941.090 -19.840 2942.270 ;
        RECT -19.420 2941.090 -18.240 2942.270 ;
        RECT -21.020 2939.490 -19.840 2940.670 ;
        RECT -19.420 2939.490 -18.240 2940.670 ;
        RECT -21.020 2761.090 -19.840 2762.270 ;
        RECT -19.420 2761.090 -18.240 2762.270 ;
        RECT -21.020 2759.490 -19.840 2760.670 ;
        RECT -19.420 2759.490 -18.240 2760.670 ;
        RECT -21.020 2581.090 -19.840 2582.270 ;
        RECT -19.420 2581.090 -18.240 2582.270 ;
        RECT -21.020 2579.490 -19.840 2580.670 ;
        RECT -19.420 2579.490 -18.240 2580.670 ;
        RECT -21.020 2401.090 -19.840 2402.270 ;
        RECT -19.420 2401.090 -18.240 2402.270 ;
        RECT -21.020 2399.490 -19.840 2400.670 ;
        RECT -19.420 2399.490 -18.240 2400.670 ;
        RECT -21.020 2221.090 -19.840 2222.270 ;
        RECT -19.420 2221.090 -18.240 2222.270 ;
        RECT -21.020 2219.490 -19.840 2220.670 ;
        RECT -19.420 2219.490 -18.240 2220.670 ;
        RECT -21.020 2041.090 -19.840 2042.270 ;
        RECT -19.420 2041.090 -18.240 2042.270 ;
        RECT -21.020 2039.490 -19.840 2040.670 ;
        RECT -19.420 2039.490 -18.240 2040.670 ;
        RECT -21.020 1861.090 -19.840 1862.270 ;
        RECT -19.420 1861.090 -18.240 1862.270 ;
        RECT -21.020 1859.490 -19.840 1860.670 ;
        RECT -19.420 1859.490 -18.240 1860.670 ;
        RECT -21.020 1681.090 -19.840 1682.270 ;
        RECT -19.420 1681.090 -18.240 1682.270 ;
        RECT -21.020 1679.490 -19.840 1680.670 ;
        RECT -19.420 1679.490 -18.240 1680.670 ;
        RECT -21.020 1501.090 -19.840 1502.270 ;
        RECT -19.420 1501.090 -18.240 1502.270 ;
        RECT -21.020 1499.490 -19.840 1500.670 ;
        RECT -19.420 1499.490 -18.240 1500.670 ;
        RECT -21.020 1321.090 -19.840 1322.270 ;
        RECT -19.420 1321.090 -18.240 1322.270 ;
        RECT -21.020 1319.490 -19.840 1320.670 ;
        RECT -19.420 1319.490 -18.240 1320.670 ;
        RECT -21.020 1141.090 -19.840 1142.270 ;
        RECT -19.420 1141.090 -18.240 1142.270 ;
        RECT -21.020 1139.490 -19.840 1140.670 ;
        RECT -19.420 1139.490 -18.240 1140.670 ;
        RECT -21.020 961.090 -19.840 962.270 ;
        RECT -19.420 961.090 -18.240 962.270 ;
        RECT -21.020 959.490 -19.840 960.670 ;
        RECT -19.420 959.490 -18.240 960.670 ;
        RECT -21.020 781.090 -19.840 782.270 ;
        RECT -19.420 781.090 -18.240 782.270 ;
        RECT -21.020 779.490 -19.840 780.670 ;
        RECT -19.420 779.490 -18.240 780.670 ;
        RECT -21.020 601.090 -19.840 602.270 ;
        RECT -19.420 601.090 -18.240 602.270 ;
        RECT -21.020 599.490 -19.840 600.670 ;
        RECT -19.420 599.490 -18.240 600.670 ;
        RECT -21.020 421.090 -19.840 422.270 ;
        RECT -19.420 421.090 -18.240 422.270 ;
        RECT -21.020 419.490 -19.840 420.670 ;
        RECT -19.420 419.490 -18.240 420.670 ;
        RECT -21.020 241.090 -19.840 242.270 ;
        RECT -19.420 241.090 -18.240 242.270 ;
        RECT -21.020 239.490 -19.840 240.670 ;
        RECT -19.420 239.490 -18.240 240.670 ;
        RECT -21.020 61.090 -19.840 62.270 ;
        RECT -19.420 61.090 -18.240 62.270 ;
        RECT -21.020 59.490 -19.840 60.670 ;
        RECT -19.420 59.490 -18.240 60.670 ;
        RECT -21.020 -14.060 -19.840 -12.880 ;
        RECT -19.420 -14.060 -18.240 -12.880 ;
        RECT -21.020 -15.660 -19.840 -14.480 ;
        RECT -19.420 -15.660 -18.240 -14.480 ;
        RECT 54.130 3534.160 55.310 3535.340 ;
        RECT 55.730 3534.160 56.910 3535.340 ;
        RECT 54.130 3532.560 55.310 3533.740 ;
        RECT 55.730 3532.560 56.910 3533.740 ;
        RECT 54.130 3481.090 55.310 3482.270 ;
        RECT 55.730 3481.090 56.910 3482.270 ;
        RECT 54.130 3479.490 55.310 3480.670 ;
        RECT 55.730 3479.490 56.910 3480.670 ;
        RECT 54.130 3301.090 55.310 3302.270 ;
        RECT 55.730 3301.090 56.910 3302.270 ;
        RECT 54.130 3299.490 55.310 3300.670 ;
        RECT 55.730 3299.490 56.910 3300.670 ;
        RECT 54.130 3121.090 55.310 3122.270 ;
        RECT 55.730 3121.090 56.910 3122.270 ;
        RECT 54.130 3119.490 55.310 3120.670 ;
        RECT 55.730 3119.490 56.910 3120.670 ;
        RECT 54.130 2941.090 55.310 2942.270 ;
        RECT 55.730 2941.090 56.910 2942.270 ;
        RECT 54.130 2939.490 55.310 2940.670 ;
        RECT 55.730 2939.490 56.910 2940.670 ;
        RECT 54.130 2761.090 55.310 2762.270 ;
        RECT 55.730 2761.090 56.910 2762.270 ;
        RECT 54.130 2759.490 55.310 2760.670 ;
        RECT 55.730 2759.490 56.910 2760.670 ;
        RECT 54.130 2581.090 55.310 2582.270 ;
        RECT 55.730 2581.090 56.910 2582.270 ;
        RECT 54.130 2579.490 55.310 2580.670 ;
        RECT 55.730 2579.490 56.910 2580.670 ;
        RECT 54.130 2401.090 55.310 2402.270 ;
        RECT 55.730 2401.090 56.910 2402.270 ;
        RECT 54.130 2399.490 55.310 2400.670 ;
        RECT 55.730 2399.490 56.910 2400.670 ;
        RECT 54.130 2221.090 55.310 2222.270 ;
        RECT 55.730 2221.090 56.910 2222.270 ;
        RECT 54.130 2219.490 55.310 2220.670 ;
        RECT 55.730 2219.490 56.910 2220.670 ;
        RECT 54.130 2041.090 55.310 2042.270 ;
        RECT 55.730 2041.090 56.910 2042.270 ;
        RECT 54.130 2039.490 55.310 2040.670 ;
        RECT 55.730 2039.490 56.910 2040.670 ;
        RECT 54.130 1861.090 55.310 1862.270 ;
        RECT 55.730 1861.090 56.910 1862.270 ;
        RECT 54.130 1859.490 55.310 1860.670 ;
        RECT 55.730 1859.490 56.910 1860.670 ;
        RECT 54.130 1681.090 55.310 1682.270 ;
        RECT 55.730 1681.090 56.910 1682.270 ;
        RECT 54.130 1679.490 55.310 1680.670 ;
        RECT 55.730 1679.490 56.910 1680.670 ;
        RECT 54.130 1501.090 55.310 1502.270 ;
        RECT 55.730 1501.090 56.910 1502.270 ;
        RECT 54.130 1499.490 55.310 1500.670 ;
        RECT 55.730 1499.490 56.910 1500.670 ;
        RECT 54.130 1321.090 55.310 1322.270 ;
        RECT 55.730 1321.090 56.910 1322.270 ;
        RECT 54.130 1319.490 55.310 1320.670 ;
        RECT 55.730 1319.490 56.910 1320.670 ;
        RECT 54.130 1141.090 55.310 1142.270 ;
        RECT 55.730 1141.090 56.910 1142.270 ;
        RECT 54.130 1139.490 55.310 1140.670 ;
        RECT 55.730 1139.490 56.910 1140.670 ;
        RECT 54.130 961.090 55.310 962.270 ;
        RECT 55.730 961.090 56.910 962.270 ;
        RECT 54.130 959.490 55.310 960.670 ;
        RECT 55.730 959.490 56.910 960.670 ;
        RECT 54.130 781.090 55.310 782.270 ;
        RECT 55.730 781.090 56.910 782.270 ;
        RECT 54.130 779.490 55.310 780.670 ;
        RECT 55.730 779.490 56.910 780.670 ;
        RECT 54.130 601.090 55.310 602.270 ;
        RECT 55.730 601.090 56.910 602.270 ;
        RECT 54.130 599.490 55.310 600.670 ;
        RECT 55.730 599.490 56.910 600.670 ;
        RECT 54.130 421.090 55.310 422.270 ;
        RECT 55.730 421.090 56.910 422.270 ;
        RECT 54.130 419.490 55.310 420.670 ;
        RECT 55.730 419.490 56.910 420.670 ;
        RECT 54.130 241.090 55.310 242.270 ;
        RECT 55.730 241.090 56.910 242.270 ;
        RECT 54.130 239.490 55.310 240.670 ;
        RECT 55.730 239.490 56.910 240.670 ;
        RECT 54.130 61.090 55.310 62.270 ;
        RECT 55.730 61.090 56.910 62.270 ;
        RECT 54.130 59.490 55.310 60.670 ;
        RECT 55.730 59.490 56.910 60.670 ;
        RECT 54.130 -14.060 55.310 -12.880 ;
        RECT 55.730 -14.060 56.910 -12.880 ;
        RECT 54.130 -15.660 55.310 -14.480 ;
        RECT 55.730 -15.660 56.910 -14.480 ;
        RECT 234.130 3534.160 235.310 3535.340 ;
        RECT 235.730 3534.160 236.910 3535.340 ;
        RECT 234.130 3532.560 235.310 3533.740 ;
        RECT 235.730 3532.560 236.910 3533.740 ;
        RECT 234.130 3481.090 235.310 3482.270 ;
        RECT 235.730 3481.090 236.910 3482.270 ;
        RECT 234.130 3479.490 235.310 3480.670 ;
        RECT 235.730 3479.490 236.910 3480.670 ;
        RECT 234.130 3301.090 235.310 3302.270 ;
        RECT 235.730 3301.090 236.910 3302.270 ;
        RECT 234.130 3299.490 235.310 3300.670 ;
        RECT 235.730 3299.490 236.910 3300.670 ;
        RECT 234.130 3121.090 235.310 3122.270 ;
        RECT 235.730 3121.090 236.910 3122.270 ;
        RECT 234.130 3119.490 235.310 3120.670 ;
        RECT 235.730 3119.490 236.910 3120.670 ;
        RECT 234.130 2941.090 235.310 2942.270 ;
        RECT 235.730 2941.090 236.910 2942.270 ;
        RECT 234.130 2939.490 235.310 2940.670 ;
        RECT 235.730 2939.490 236.910 2940.670 ;
        RECT 234.130 2761.090 235.310 2762.270 ;
        RECT 235.730 2761.090 236.910 2762.270 ;
        RECT 234.130 2759.490 235.310 2760.670 ;
        RECT 235.730 2759.490 236.910 2760.670 ;
        RECT 234.130 2581.090 235.310 2582.270 ;
        RECT 235.730 2581.090 236.910 2582.270 ;
        RECT 234.130 2579.490 235.310 2580.670 ;
        RECT 235.730 2579.490 236.910 2580.670 ;
        RECT 234.130 2401.090 235.310 2402.270 ;
        RECT 235.730 2401.090 236.910 2402.270 ;
        RECT 234.130 2399.490 235.310 2400.670 ;
        RECT 235.730 2399.490 236.910 2400.670 ;
        RECT 234.130 2221.090 235.310 2222.270 ;
        RECT 235.730 2221.090 236.910 2222.270 ;
        RECT 234.130 2219.490 235.310 2220.670 ;
        RECT 235.730 2219.490 236.910 2220.670 ;
        RECT 234.130 2041.090 235.310 2042.270 ;
        RECT 235.730 2041.090 236.910 2042.270 ;
        RECT 234.130 2039.490 235.310 2040.670 ;
        RECT 235.730 2039.490 236.910 2040.670 ;
        RECT 234.130 1861.090 235.310 1862.270 ;
        RECT 235.730 1861.090 236.910 1862.270 ;
        RECT 234.130 1859.490 235.310 1860.670 ;
        RECT 235.730 1859.490 236.910 1860.670 ;
        RECT 234.130 1681.090 235.310 1682.270 ;
        RECT 235.730 1681.090 236.910 1682.270 ;
        RECT 234.130 1679.490 235.310 1680.670 ;
        RECT 235.730 1679.490 236.910 1680.670 ;
        RECT 234.130 1501.090 235.310 1502.270 ;
        RECT 235.730 1501.090 236.910 1502.270 ;
        RECT 234.130 1499.490 235.310 1500.670 ;
        RECT 235.730 1499.490 236.910 1500.670 ;
        RECT 234.130 1321.090 235.310 1322.270 ;
        RECT 235.730 1321.090 236.910 1322.270 ;
        RECT 234.130 1319.490 235.310 1320.670 ;
        RECT 235.730 1319.490 236.910 1320.670 ;
        RECT 234.130 1141.090 235.310 1142.270 ;
        RECT 235.730 1141.090 236.910 1142.270 ;
        RECT 234.130 1139.490 235.310 1140.670 ;
        RECT 235.730 1139.490 236.910 1140.670 ;
        RECT 234.130 961.090 235.310 962.270 ;
        RECT 235.730 961.090 236.910 962.270 ;
        RECT 234.130 959.490 235.310 960.670 ;
        RECT 235.730 959.490 236.910 960.670 ;
        RECT 234.130 781.090 235.310 782.270 ;
        RECT 235.730 781.090 236.910 782.270 ;
        RECT 234.130 779.490 235.310 780.670 ;
        RECT 235.730 779.490 236.910 780.670 ;
        RECT 414.130 3534.160 415.310 3535.340 ;
        RECT 415.730 3534.160 416.910 3535.340 ;
        RECT 414.130 3532.560 415.310 3533.740 ;
        RECT 415.730 3532.560 416.910 3533.740 ;
        RECT 414.130 3481.090 415.310 3482.270 ;
        RECT 415.730 3481.090 416.910 3482.270 ;
        RECT 414.130 3479.490 415.310 3480.670 ;
        RECT 415.730 3479.490 416.910 3480.670 ;
        RECT 414.130 3301.090 415.310 3302.270 ;
        RECT 415.730 3301.090 416.910 3302.270 ;
        RECT 414.130 3299.490 415.310 3300.670 ;
        RECT 415.730 3299.490 416.910 3300.670 ;
        RECT 414.130 3121.090 415.310 3122.270 ;
        RECT 415.730 3121.090 416.910 3122.270 ;
        RECT 414.130 3119.490 415.310 3120.670 ;
        RECT 415.730 3119.490 416.910 3120.670 ;
        RECT 414.130 2941.090 415.310 2942.270 ;
        RECT 415.730 2941.090 416.910 2942.270 ;
        RECT 414.130 2939.490 415.310 2940.670 ;
        RECT 415.730 2939.490 416.910 2940.670 ;
        RECT 414.130 2761.090 415.310 2762.270 ;
        RECT 415.730 2761.090 416.910 2762.270 ;
        RECT 414.130 2759.490 415.310 2760.670 ;
        RECT 415.730 2759.490 416.910 2760.670 ;
        RECT 414.130 2581.090 415.310 2582.270 ;
        RECT 415.730 2581.090 416.910 2582.270 ;
        RECT 414.130 2579.490 415.310 2580.670 ;
        RECT 415.730 2579.490 416.910 2580.670 ;
        RECT 414.130 2401.090 415.310 2402.270 ;
        RECT 415.730 2401.090 416.910 2402.270 ;
        RECT 414.130 2399.490 415.310 2400.670 ;
        RECT 415.730 2399.490 416.910 2400.670 ;
        RECT 414.130 2221.090 415.310 2222.270 ;
        RECT 415.730 2221.090 416.910 2222.270 ;
        RECT 414.130 2219.490 415.310 2220.670 ;
        RECT 415.730 2219.490 416.910 2220.670 ;
        RECT 414.130 2041.090 415.310 2042.270 ;
        RECT 415.730 2041.090 416.910 2042.270 ;
        RECT 414.130 2039.490 415.310 2040.670 ;
        RECT 415.730 2039.490 416.910 2040.670 ;
        RECT 414.130 1861.090 415.310 1862.270 ;
        RECT 415.730 1861.090 416.910 1862.270 ;
        RECT 414.130 1859.490 415.310 1860.670 ;
        RECT 415.730 1859.490 416.910 1860.670 ;
        RECT 414.130 1681.090 415.310 1682.270 ;
        RECT 415.730 1681.090 416.910 1682.270 ;
        RECT 414.130 1679.490 415.310 1680.670 ;
        RECT 415.730 1679.490 416.910 1680.670 ;
        RECT 414.130 1501.090 415.310 1502.270 ;
        RECT 415.730 1501.090 416.910 1502.270 ;
        RECT 414.130 1499.490 415.310 1500.670 ;
        RECT 415.730 1499.490 416.910 1500.670 ;
        RECT 414.130 1321.090 415.310 1322.270 ;
        RECT 415.730 1321.090 416.910 1322.270 ;
        RECT 414.130 1319.490 415.310 1320.670 ;
        RECT 415.730 1319.490 416.910 1320.670 ;
        RECT 414.130 1141.090 415.310 1142.270 ;
        RECT 415.730 1141.090 416.910 1142.270 ;
        RECT 414.130 1139.490 415.310 1140.670 ;
        RECT 415.730 1139.490 416.910 1140.670 ;
        RECT 414.130 961.090 415.310 962.270 ;
        RECT 415.730 961.090 416.910 962.270 ;
        RECT 414.130 959.490 415.310 960.670 ;
        RECT 415.730 959.490 416.910 960.670 ;
        RECT 414.130 781.090 415.310 782.270 ;
        RECT 415.730 781.090 416.910 782.270 ;
        RECT 414.130 779.490 415.310 780.670 ;
        RECT 415.730 779.490 416.910 780.670 ;
        RECT 594.130 3534.160 595.310 3535.340 ;
        RECT 595.730 3534.160 596.910 3535.340 ;
        RECT 594.130 3532.560 595.310 3533.740 ;
        RECT 595.730 3532.560 596.910 3533.740 ;
        RECT 594.130 3481.090 595.310 3482.270 ;
        RECT 595.730 3481.090 596.910 3482.270 ;
        RECT 594.130 3479.490 595.310 3480.670 ;
        RECT 595.730 3479.490 596.910 3480.670 ;
        RECT 594.130 3301.090 595.310 3302.270 ;
        RECT 595.730 3301.090 596.910 3302.270 ;
        RECT 594.130 3299.490 595.310 3300.670 ;
        RECT 595.730 3299.490 596.910 3300.670 ;
        RECT 594.130 3121.090 595.310 3122.270 ;
        RECT 595.730 3121.090 596.910 3122.270 ;
        RECT 594.130 3119.490 595.310 3120.670 ;
        RECT 595.730 3119.490 596.910 3120.670 ;
        RECT 594.130 2941.090 595.310 2942.270 ;
        RECT 595.730 2941.090 596.910 2942.270 ;
        RECT 594.130 2939.490 595.310 2940.670 ;
        RECT 595.730 2939.490 596.910 2940.670 ;
        RECT 594.130 2761.090 595.310 2762.270 ;
        RECT 595.730 2761.090 596.910 2762.270 ;
        RECT 594.130 2759.490 595.310 2760.670 ;
        RECT 595.730 2759.490 596.910 2760.670 ;
        RECT 594.130 2581.090 595.310 2582.270 ;
        RECT 595.730 2581.090 596.910 2582.270 ;
        RECT 594.130 2579.490 595.310 2580.670 ;
        RECT 595.730 2579.490 596.910 2580.670 ;
        RECT 594.130 2401.090 595.310 2402.270 ;
        RECT 595.730 2401.090 596.910 2402.270 ;
        RECT 594.130 2399.490 595.310 2400.670 ;
        RECT 595.730 2399.490 596.910 2400.670 ;
        RECT 594.130 2221.090 595.310 2222.270 ;
        RECT 595.730 2221.090 596.910 2222.270 ;
        RECT 594.130 2219.490 595.310 2220.670 ;
        RECT 595.730 2219.490 596.910 2220.670 ;
        RECT 594.130 2041.090 595.310 2042.270 ;
        RECT 595.730 2041.090 596.910 2042.270 ;
        RECT 594.130 2039.490 595.310 2040.670 ;
        RECT 595.730 2039.490 596.910 2040.670 ;
        RECT 594.130 1861.090 595.310 1862.270 ;
        RECT 595.730 1861.090 596.910 1862.270 ;
        RECT 594.130 1859.490 595.310 1860.670 ;
        RECT 595.730 1859.490 596.910 1860.670 ;
        RECT 594.130 1681.090 595.310 1682.270 ;
        RECT 595.730 1681.090 596.910 1682.270 ;
        RECT 594.130 1679.490 595.310 1680.670 ;
        RECT 595.730 1679.490 596.910 1680.670 ;
        RECT 594.130 1501.090 595.310 1502.270 ;
        RECT 595.730 1501.090 596.910 1502.270 ;
        RECT 594.130 1499.490 595.310 1500.670 ;
        RECT 595.730 1499.490 596.910 1500.670 ;
        RECT 594.130 1321.090 595.310 1322.270 ;
        RECT 595.730 1321.090 596.910 1322.270 ;
        RECT 594.130 1319.490 595.310 1320.670 ;
        RECT 595.730 1319.490 596.910 1320.670 ;
        RECT 594.130 1141.090 595.310 1142.270 ;
        RECT 595.730 1141.090 596.910 1142.270 ;
        RECT 594.130 1139.490 595.310 1140.670 ;
        RECT 595.730 1139.490 596.910 1140.670 ;
        RECT 594.130 961.090 595.310 962.270 ;
        RECT 595.730 961.090 596.910 962.270 ;
        RECT 594.130 959.490 595.310 960.670 ;
        RECT 595.730 959.490 596.910 960.670 ;
        RECT 594.130 781.090 595.310 782.270 ;
        RECT 595.730 781.090 596.910 782.270 ;
        RECT 594.130 779.490 595.310 780.670 ;
        RECT 595.730 779.490 596.910 780.670 ;
        RECT 774.130 3534.160 775.310 3535.340 ;
        RECT 775.730 3534.160 776.910 3535.340 ;
        RECT 774.130 3532.560 775.310 3533.740 ;
        RECT 775.730 3532.560 776.910 3533.740 ;
        RECT 774.130 3481.090 775.310 3482.270 ;
        RECT 775.730 3481.090 776.910 3482.270 ;
        RECT 774.130 3479.490 775.310 3480.670 ;
        RECT 775.730 3479.490 776.910 3480.670 ;
        RECT 774.130 3301.090 775.310 3302.270 ;
        RECT 775.730 3301.090 776.910 3302.270 ;
        RECT 774.130 3299.490 775.310 3300.670 ;
        RECT 775.730 3299.490 776.910 3300.670 ;
        RECT 774.130 3121.090 775.310 3122.270 ;
        RECT 775.730 3121.090 776.910 3122.270 ;
        RECT 774.130 3119.490 775.310 3120.670 ;
        RECT 775.730 3119.490 776.910 3120.670 ;
        RECT 774.130 2941.090 775.310 2942.270 ;
        RECT 775.730 2941.090 776.910 2942.270 ;
        RECT 774.130 2939.490 775.310 2940.670 ;
        RECT 775.730 2939.490 776.910 2940.670 ;
        RECT 774.130 2761.090 775.310 2762.270 ;
        RECT 775.730 2761.090 776.910 2762.270 ;
        RECT 774.130 2759.490 775.310 2760.670 ;
        RECT 775.730 2759.490 776.910 2760.670 ;
        RECT 774.130 2581.090 775.310 2582.270 ;
        RECT 775.730 2581.090 776.910 2582.270 ;
        RECT 774.130 2579.490 775.310 2580.670 ;
        RECT 775.730 2579.490 776.910 2580.670 ;
        RECT 774.130 2401.090 775.310 2402.270 ;
        RECT 775.730 2401.090 776.910 2402.270 ;
        RECT 774.130 2399.490 775.310 2400.670 ;
        RECT 775.730 2399.490 776.910 2400.670 ;
        RECT 774.130 2221.090 775.310 2222.270 ;
        RECT 775.730 2221.090 776.910 2222.270 ;
        RECT 774.130 2219.490 775.310 2220.670 ;
        RECT 775.730 2219.490 776.910 2220.670 ;
        RECT 774.130 2041.090 775.310 2042.270 ;
        RECT 775.730 2041.090 776.910 2042.270 ;
        RECT 774.130 2039.490 775.310 2040.670 ;
        RECT 775.730 2039.490 776.910 2040.670 ;
        RECT 774.130 1861.090 775.310 1862.270 ;
        RECT 775.730 1861.090 776.910 1862.270 ;
        RECT 774.130 1859.490 775.310 1860.670 ;
        RECT 775.730 1859.490 776.910 1860.670 ;
        RECT 774.130 1681.090 775.310 1682.270 ;
        RECT 775.730 1681.090 776.910 1682.270 ;
        RECT 774.130 1679.490 775.310 1680.670 ;
        RECT 775.730 1679.490 776.910 1680.670 ;
        RECT 774.130 1501.090 775.310 1502.270 ;
        RECT 775.730 1501.090 776.910 1502.270 ;
        RECT 774.130 1499.490 775.310 1500.670 ;
        RECT 775.730 1499.490 776.910 1500.670 ;
        RECT 774.130 1321.090 775.310 1322.270 ;
        RECT 775.730 1321.090 776.910 1322.270 ;
        RECT 774.130 1319.490 775.310 1320.670 ;
        RECT 775.730 1319.490 776.910 1320.670 ;
        RECT 774.130 1141.090 775.310 1142.270 ;
        RECT 775.730 1141.090 776.910 1142.270 ;
        RECT 774.130 1139.490 775.310 1140.670 ;
        RECT 775.730 1139.490 776.910 1140.670 ;
        RECT 774.130 961.090 775.310 962.270 ;
        RECT 775.730 961.090 776.910 962.270 ;
        RECT 774.130 959.490 775.310 960.670 ;
        RECT 775.730 959.490 776.910 960.670 ;
        RECT 774.130 781.090 775.310 782.270 ;
        RECT 775.730 781.090 776.910 782.270 ;
        RECT 774.130 779.490 775.310 780.670 ;
        RECT 775.730 779.490 776.910 780.670 ;
        RECT 234.130 601.090 235.310 602.270 ;
        RECT 235.730 601.090 236.910 602.270 ;
        RECT 234.130 599.490 235.310 600.670 ;
        RECT 235.730 599.490 236.910 600.670 ;
        RECT 774.130 601.090 775.310 602.270 ;
        RECT 775.730 601.090 776.910 602.270 ;
        RECT 774.130 599.490 775.310 600.670 ;
        RECT 775.730 599.490 776.910 600.670 ;
        RECT 234.130 421.090 235.310 422.270 ;
        RECT 235.730 421.090 236.910 422.270 ;
        RECT 234.130 419.490 235.310 420.670 ;
        RECT 235.730 419.490 236.910 420.670 ;
        RECT 234.130 241.090 235.310 242.270 ;
        RECT 235.730 241.090 236.910 242.270 ;
        RECT 234.130 239.490 235.310 240.670 ;
        RECT 235.730 239.490 236.910 240.670 ;
        RECT 234.130 61.090 235.310 62.270 ;
        RECT 235.730 61.090 236.910 62.270 ;
        RECT 234.130 59.490 235.310 60.670 ;
        RECT 235.730 59.490 236.910 60.670 ;
        RECT 234.130 -14.060 235.310 -12.880 ;
        RECT 235.730 -14.060 236.910 -12.880 ;
        RECT 234.130 -15.660 235.310 -14.480 ;
        RECT 235.730 -15.660 236.910 -14.480 ;
        RECT 414.130 421.090 415.310 422.270 ;
        RECT 415.730 421.090 416.910 422.270 ;
        RECT 414.130 419.490 415.310 420.670 ;
        RECT 415.730 419.490 416.910 420.670 ;
        RECT 414.130 241.090 415.310 242.270 ;
        RECT 415.730 241.090 416.910 242.270 ;
        RECT 414.130 239.490 415.310 240.670 ;
        RECT 415.730 239.490 416.910 240.670 ;
        RECT 414.130 61.090 415.310 62.270 ;
        RECT 415.730 61.090 416.910 62.270 ;
        RECT 414.130 59.490 415.310 60.670 ;
        RECT 415.730 59.490 416.910 60.670 ;
        RECT 414.130 -14.060 415.310 -12.880 ;
        RECT 415.730 -14.060 416.910 -12.880 ;
        RECT 414.130 -15.660 415.310 -14.480 ;
        RECT 415.730 -15.660 416.910 -14.480 ;
        RECT 594.130 421.090 595.310 422.270 ;
        RECT 595.730 421.090 596.910 422.270 ;
        RECT 594.130 419.490 595.310 420.670 ;
        RECT 595.730 419.490 596.910 420.670 ;
        RECT 594.130 241.090 595.310 242.270 ;
        RECT 595.730 241.090 596.910 242.270 ;
        RECT 594.130 239.490 595.310 240.670 ;
        RECT 595.730 239.490 596.910 240.670 ;
        RECT 594.130 61.090 595.310 62.270 ;
        RECT 595.730 61.090 596.910 62.270 ;
        RECT 594.130 59.490 595.310 60.670 ;
        RECT 595.730 59.490 596.910 60.670 ;
        RECT 594.130 -14.060 595.310 -12.880 ;
        RECT 595.730 -14.060 596.910 -12.880 ;
        RECT 594.130 -15.660 595.310 -14.480 ;
        RECT 595.730 -15.660 596.910 -14.480 ;
        RECT 774.130 421.090 775.310 422.270 ;
        RECT 775.730 421.090 776.910 422.270 ;
        RECT 774.130 419.490 775.310 420.670 ;
        RECT 775.730 419.490 776.910 420.670 ;
        RECT 774.130 241.090 775.310 242.270 ;
        RECT 775.730 241.090 776.910 242.270 ;
        RECT 774.130 239.490 775.310 240.670 ;
        RECT 775.730 239.490 776.910 240.670 ;
        RECT 774.130 61.090 775.310 62.270 ;
        RECT 775.730 61.090 776.910 62.270 ;
        RECT 774.130 59.490 775.310 60.670 ;
        RECT 775.730 59.490 776.910 60.670 ;
        RECT 774.130 -14.060 775.310 -12.880 ;
        RECT 775.730 -14.060 776.910 -12.880 ;
        RECT 774.130 -15.660 775.310 -14.480 ;
        RECT 775.730 -15.660 776.910 -14.480 ;
        RECT 954.130 3534.160 955.310 3535.340 ;
        RECT 955.730 3534.160 956.910 3535.340 ;
        RECT 954.130 3532.560 955.310 3533.740 ;
        RECT 955.730 3532.560 956.910 3533.740 ;
        RECT 954.130 3481.090 955.310 3482.270 ;
        RECT 955.730 3481.090 956.910 3482.270 ;
        RECT 954.130 3479.490 955.310 3480.670 ;
        RECT 955.730 3479.490 956.910 3480.670 ;
        RECT 954.130 3301.090 955.310 3302.270 ;
        RECT 955.730 3301.090 956.910 3302.270 ;
        RECT 954.130 3299.490 955.310 3300.670 ;
        RECT 955.730 3299.490 956.910 3300.670 ;
        RECT 954.130 3121.090 955.310 3122.270 ;
        RECT 955.730 3121.090 956.910 3122.270 ;
        RECT 954.130 3119.490 955.310 3120.670 ;
        RECT 955.730 3119.490 956.910 3120.670 ;
        RECT 954.130 2941.090 955.310 2942.270 ;
        RECT 955.730 2941.090 956.910 2942.270 ;
        RECT 954.130 2939.490 955.310 2940.670 ;
        RECT 955.730 2939.490 956.910 2940.670 ;
        RECT 954.130 2761.090 955.310 2762.270 ;
        RECT 955.730 2761.090 956.910 2762.270 ;
        RECT 954.130 2759.490 955.310 2760.670 ;
        RECT 955.730 2759.490 956.910 2760.670 ;
        RECT 954.130 2581.090 955.310 2582.270 ;
        RECT 955.730 2581.090 956.910 2582.270 ;
        RECT 954.130 2579.490 955.310 2580.670 ;
        RECT 955.730 2579.490 956.910 2580.670 ;
        RECT 954.130 2401.090 955.310 2402.270 ;
        RECT 955.730 2401.090 956.910 2402.270 ;
        RECT 954.130 2399.490 955.310 2400.670 ;
        RECT 955.730 2399.490 956.910 2400.670 ;
        RECT 954.130 2221.090 955.310 2222.270 ;
        RECT 955.730 2221.090 956.910 2222.270 ;
        RECT 954.130 2219.490 955.310 2220.670 ;
        RECT 955.730 2219.490 956.910 2220.670 ;
        RECT 954.130 2041.090 955.310 2042.270 ;
        RECT 955.730 2041.090 956.910 2042.270 ;
        RECT 954.130 2039.490 955.310 2040.670 ;
        RECT 955.730 2039.490 956.910 2040.670 ;
        RECT 954.130 1861.090 955.310 1862.270 ;
        RECT 955.730 1861.090 956.910 1862.270 ;
        RECT 954.130 1859.490 955.310 1860.670 ;
        RECT 955.730 1859.490 956.910 1860.670 ;
        RECT 954.130 1681.090 955.310 1682.270 ;
        RECT 955.730 1681.090 956.910 1682.270 ;
        RECT 954.130 1679.490 955.310 1680.670 ;
        RECT 955.730 1679.490 956.910 1680.670 ;
        RECT 954.130 1501.090 955.310 1502.270 ;
        RECT 955.730 1501.090 956.910 1502.270 ;
        RECT 954.130 1499.490 955.310 1500.670 ;
        RECT 955.730 1499.490 956.910 1500.670 ;
        RECT 954.130 1321.090 955.310 1322.270 ;
        RECT 955.730 1321.090 956.910 1322.270 ;
        RECT 954.130 1319.490 955.310 1320.670 ;
        RECT 955.730 1319.490 956.910 1320.670 ;
        RECT 954.130 1141.090 955.310 1142.270 ;
        RECT 955.730 1141.090 956.910 1142.270 ;
        RECT 954.130 1139.490 955.310 1140.670 ;
        RECT 955.730 1139.490 956.910 1140.670 ;
        RECT 954.130 961.090 955.310 962.270 ;
        RECT 955.730 961.090 956.910 962.270 ;
        RECT 954.130 959.490 955.310 960.670 ;
        RECT 955.730 959.490 956.910 960.670 ;
        RECT 954.130 781.090 955.310 782.270 ;
        RECT 955.730 781.090 956.910 782.270 ;
        RECT 954.130 779.490 955.310 780.670 ;
        RECT 955.730 779.490 956.910 780.670 ;
        RECT 954.130 601.090 955.310 602.270 ;
        RECT 955.730 601.090 956.910 602.270 ;
        RECT 954.130 599.490 955.310 600.670 ;
        RECT 955.730 599.490 956.910 600.670 ;
        RECT 954.130 421.090 955.310 422.270 ;
        RECT 955.730 421.090 956.910 422.270 ;
        RECT 954.130 419.490 955.310 420.670 ;
        RECT 955.730 419.490 956.910 420.670 ;
        RECT 954.130 241.090 955.310 242.270 ;
        RECT 955.730 241.090 956.910 242.270 ;
        RECT 954.130 239.490 955.310 240.670 ;
        RECT 955.730 239.490 956.910 240.670 ;
        RECT 954.130 61.090 955.310 62.270 ;
        RECT 955.730 61.090 956.910 62.270 ;
        RECT 954.130 59.490 955.310 60.670 ;
        RECT 955.730 59.490 956.910 60.670 ;
        RECT 954.130 -14.060 955.310 -12.880 ;
        RECT 955.730 -14.060 956.910 -12.880 ;
        RECT 954.130 -15.660 955.310 -14.480 ;
        RECT 955.730 -15.660 956.910 -14.480 ;
        RECT 1134.130 3534.160 1135.310 3535.340 ;
        RECT 1135.730 3534.160 1136.910 3535.340 ;
        RECT 1134.130 3532.560 1135.310 3533.740 ;
        RECT 1135.730 3532.560 1136.910 3533.740 ;
        RECT 1134.130 3481.090 1135.310 3482.270 ;
        RECT 1135.730 3481.090 1136.910 3482.270 ;
        RECT 1134.130 3479.490 1135.310 3480.670 ;
        RECT 1135.730 3479.490 1136.910 3480.670 ;
        RECT 1134.130 3301.090 1135.310 3302.270 ;
        RECT 1135.730 3301.090 1136.910 3302.270 ;
        RECT 1134.130 3299.490 1135.310 3300.670 ;
        RECT 1135.730 3299.490 1136.910 3300.670 ;
        RECT 1134.130 3121.090 1135.310 3122.270 ;
        RECT 1135.730 3121.090 1136.910 3122.270 ;
        RECT 1134.130 3119.490 1135.310 3120.670 ;
        RECT 1135.730 3119.490 1136.910 3120.670 ;
        RECT 1134.130 2941.090 1135.310 2942.270 ;
        RECT 1135.730 2941.090 1136.910 2942.270 ;
        RECT 1134.130 2939.490 1135.310 2940.670 ;
        RECT 1135.730 2939.490 1136.910 2940.670 ;
        RECT 1134.130 2761.090 1135.310 2762.270 ;
        RECT 1135.730 2761.090 1136.910 2762.270 ;
        RECT 1134.130 2759.490 1135.310 2760.670 ;
        RECT 1135.730 2759.490 1136.910 2760.670 ;
        RECT 1134.130 2581.090 1135.310 2582.270 ;
        RECT 1135.730 2581.090 1136.910 2582.270 ;
        RECT 1134.130 2579.490 1135.310 2580.670 ;
        RECT 1135.730 2579.490 1136.910 2580.670 ;
        RECT 1134.130 2401.090 1135.310 2402.270 ;
        RECT 1135.730 2401.090 1136.910 2402.270 ;
        RECT 1134.130 2399.490 1135.310 2400.670 ;
        RECT 1135.730 2399.490 1136.910 2400.670 ;
        RECT 1134.130 2221.090 1135.310 2222.270 ;
        RECT 1135.730 2221.090 1136.910 2222.270 ;
        RECT 1134.130 2219.490 1135.310 2220.670 ;
        RECT 1135.730 2219.490 1136.910 2220.670 ;
        RECT 1134.130 2041.090 1135.310 2042.270 ;
        RECT 1135.730 2041.090 1136.910 2042.270 ;
        RECT 1134.130 2039.490 1135.310 2040.670 ;
        RECT 1135.730 2039.490 1136.910 2040.670 ;
        RECT 1134.130 1861.090 1135.310 1862.270 ;
        RECT 1135.730 1861.090 1136.910 1862.270 ;
        RECT 1134.130 1859.490 1135.310 1860.670 ;
        RECT 1135.730 1859.490 1136.910 1860.670 ;
        RECT 1134.130 1681.090 1135.310 1682.270 ;
        RECT 1135.730 1681.090 1136.910 1682.270 ;
        RECT 1134.130 1679.490 1135.310 1680.670 ;
        RECT 1135.730 1679.490 1136.910 1680.670 ;
        RECT 1134.130 1501.090 1135.310 1502.270 ;
        RECT 1135.730 1501.090 1136.910 1502.270 ;
        RECT 1134.130 1499.490 1135.310 1500.670 ;
        RECT 1135.730 1499.490 1136.910 1500.670 ;
        RECT 1134.130 1321.090 1135.310 1322.270 ;
        RECT 1135.730 1321.090 1136.910 1322.270 ;
        RECT 1134.130 1319.490 1135.310 1320.670 ;
        RECT 1135.730 1319.490 1136.910 1320.670 ;
        RECT 1134.130 1141.090 1135.310 1142.270 ;
        RECT 1135.730 1141.090 1136.910 1142.270 ;
        RECT 1134.130 1139.490 1135.310 1140.670 ;
        RECT 1135.730 1139.490 1136.910 1140.670 ;
        RECT 1134.130 961.090 1135.310 962.270 ;
        RECT 1135.730 961.090 1136.910 962.270 ;
        RECT 1134.130 959.490 1135.310 960.670 ;
        RECT 1135.730 959.490 1136.910 960.670 ;
        RECT 1134.130 781.090 1135.310 782.270 ;
        RECT 1135.730 781.090 1136.910 782.270 ;
        RECT 1134.130 779.490 1135.310 780.670 ;
        RECT 1135.730 779.490 1136.910 780.670 ;
        RECT 1134.130 601.090 1135.310 602.270 ;
        RECT 1135.730 601.090 1136.910 602.270 ;
        RECT 1134.130 599.490 1135.310 600.670 ;
        RECT 1135.730 599.490 1136.910 600.670 ;
        RECT 1134.130 421.090 1135.310 422.270 ;
        RECT 1135.730 421.090 1136.910 422.270 ;
        RECT 1134.130 419.490 1135.310 420.670 ;
        RECT 1135.730 419.490 1136.910 420.670 ;
        RECT 1134.130 241.090 1135.310 242.270 ;
        RECT 1135.730 241.090 1136.910 242.270 ;
        RECT 1134.130 239.490 1135.310 240.670 ;
        RECT 1135.730 239.490 1136.910 240.670 ;
        RECT 1134.130 61.090 1135.310 62.270 ;
        RECT 1135.730 61.090 1136.910 62.270 ;
        RECT 1134.130 59.490 1135.310 60.670 ;
        RECT 1135.730 59.490 1136.910 60.670 ;
        RECT 1134.130 -14.060 1135.310 -12.880 ;
        RECT 1135.730 -14.060 1136.910 -12.880 ;
        RECT 1134.130 -15.660 1135.310 -14.480 ;
        RECT 1135.730 -15.660 1136.910 -14.480 ;
        RECT 1314.130 3534.160 1315.310 3535.340 ;
        RECT 1315.730 3534.160 1316.910 3535.340 ;
        RECT 1314.130 3532.560 1315.310 3533.740 ;
        RECT 1315.730 3532.560 1316.910 3533.740 ;
        RECT 1314.130 3481.090 1315.310 3482.270 ;
        RECT 1315.730 3481.090 1316.910 3482.270 ;
        RECT 1314.130 3479.490 1315.310 3480.670 ;
        RECT 1315.730 3479.490 1316.910 3480.670 ;
        RECT 1314.130 3301.090 1315.310 3302.270 ;
        RECT 1315.730 3301.090 1316.910 3302.270 ;
        RECT 1314.130 3299.490 1315.310 3300.670 ;
        RECT 1315.730 3299.490 1316.910 3300.670 ;
        RECT 1314.130 3121.090 1315.310 3122.270 ;
        RECT 1315.730 3121.090 1316.910 3122.270 ;
        RECT 1314.130 3119.490 1315.310 3120.670 ;
        RECT 1315.730 3119.490 1316.910 3120.670 ;
        RECT 1314.130 2941.090 1315.310 2942.270 ;
        RECT 1315.730 2941.090 1316.910 2942.270 ;
        RECT 1314.130 2939.490 1315.310 2940.670 ;
        RECT 1315.730 2939.490 1316.910 2940.670 ;
        RECT 1314.130 2761.090 1315.310 2762.270 ;
        RECT 1315.730 2761.090 1316.910 2762.270 ;
        RECT 1314.130 2759.490 1315.310 2760.670 ;
        RECT 1315.730 2759.490 1316.910 2760.670 ;
        RECT 1314.130 2581.090 1315.310 2582.270 ;
        RECT 1315.730 2581.090 1316.910 2582.270 ;
        RECT 1314.130 2579.490 1315.310 2580.670 ;
        RECT 1315.730 2579.490 1316.910 2580.670 ;
        RECT 1314.130 2401.090 1315.310 2402.270 ;
        RECT 1315.730 2401.090 1316.910 2402.270 ;
        RECT 1314.130 2399.490 1315.310 2400.670 ;
        RECT 1315.730 2399.490 1316.910 2400.670 ;
        RECT 1314.130 2221.090 1315.310 2222.270 ;
        RECT 1315.730 2221.090 1316.910 2222.270 ;
        RECT 1314.130 2219.490 1315.310 2220.670 ;
        RECT 1315.730 2219.490 1316.910 2220.670 ;
        RECT 1314.130 2041.090 1315.310 2042.270 ;
        RECT 1315.730 2041.090 1316.910 2042.270 ;
        RECT 1314.130 2039.490 1315.310 2040.670 ;
        RECT 1315.730 2039.490 1316.910 2040.670 ;
        RECT 1314.130 1861.090 1315.310 1862.270 ;
        RECT 1315.730 1861.090 1316.910 1862.270 ;
        RECT 1314.130 1859.490 1315.310 1860.670 ;
        RECT 1315.730 1859.490 1316.910 1860.670 ;
        RECT 1314.130 1681.090 1315.310 1682.270 ;
        RECT 1315.730 1681.090 1316.910 1682.270 ;
        RECT 1314.130 1679.490 1315.310 1680.670 ;
        RECT 1315.730 1679.490 1316.910 1680.670 ;
        RECT 1314.130 1501.090 1315.310 1502.270 ;
        RECT 1315.730 1501.090 1316.910 1502.270 ;
        RECT 1314.130 1499.490 1315.310 1500.670 ;
        RECT 1315.730 1499.490 1316.910 1500.670 ;
        RECT 1314.130 1321.090 1315.310 1322.270 ;
        RECT 1315.730 1321.090 1316.910 1322.270 ;
        RECT 1314.130 1319.490 1315.310 1320.670 ;
        RECT 1315.730 1319.490 1316.910 1320.670 ;
        RECT 1314.130 1141.090 1315.310 1142.270 ;
        RECT 1315.730 1141.090 1316.910 1142.270 ;
        RECT 1314.130 1139.490 1315.310 1140.670 ;
        RECT 1315.730 1139.490 1316.910 1140.670 ;
        RECT 1314.130 961.090 1315.310 962.270 ;
        RECT 1315.730 961.090 1316.910 962.270 ;
        RECT 1314.130 959.490 1315.310 960.670 ;
        RECT 1315.730 959.490 1316.910 960.670 ;
        RECT 1314.130 781.090 1315.310 782.270 ;
        RECT 1315.730 781.090 1316.910 782.270 ;
        RECT 1314.130 779.490 1315.310 780.670 ;
        RECT 1315.730 779.490 1316.910 780.670 ;
        RECT 1314.130 601.090 1315.310 602.270 ;
        RECT 1315.730 601.090 1316.910 602.270 ;
        RECT 1314.130 599.490 1315.310 600.670 ;
        RECT 1315.730 599.490 1316.910 600.670 ;
        RECT 1314.130 421.090 1315.310 422.270 ;
        RECT 1315.730 421.090 1316.910 422.270 ;
        RECT 1314.130 419.490 1315.310 420.670 ;
        RECT 1315.730 419.490 1316.910 420.670 ;
        RECT 1314.130 241.090 1315.310 242.270 ;
        RECT 1315.730 241.090 1316.910 242.270 ;
        RECT 1314.130 239.490 1315.310 240.670 ;
        RECT 1315.730 239.490 1316.910 240.670 ;
        RECT 1314.130 61.090 1315.310 62.270 ;
        RECT 1315.730 61.090 1316.910 62.270 ;
        RECT 1314.130 59.490 1315.310 60.670 ;
        RECT 1315.730 59.490 1316.910 60.670 ;
        RECT 1314.130 -14.060 1315.310 -12.880 ;
        RECT 1315.730 -14.060 1316.910 -12.880 ;
        RECT 1314.130 -15.660 1315.310 -14.480 ;
        RECT 1315.730 -15.660 1316.910 -14.480 ;
        RECT 1494.130 3534.160 1495.310 3535.340 ;
        RECT 1495.730 3534.160 1496.910 3535.340 ;
        RECT 1494.130 3532.560 1495.310 3533.740 ;
        RECT 1495.730 3532.560 1496.910 3533.740 ;
        RECT 1494.130 3481.090 1495.310 3482.270 ;
        RECT 1495.730 3481.090 1496.910 3482.270 ;
        RECT 1494.130 3479.490 1495.310 3480.670 ;
        RECT 1495.730 3479.490 1496.910 3480.670 ;
        RECT 1494.130 3301.090 1495.310 3302.270 ;
        RECT 1495.730 3301.090 1496.910 3302.270 ;
        RECT 1494.130 3299.490 1495.310 3300.670 ;
        RECT 1495.730 3299.490 1496.910 3300.670 ;
        RECT 1494.130 3121.090 1495.310 3122.270 ;
        RECT 1495.730 3121.090 1496.910 3122.270 ;
        RECT 1494.130 3119.490 1495.310 3120.670 ;
        RECT 1495.730 3119.490 1496.910 3120.670 ;
        RECT 1494.130 2941.090 1495.310 2942.270 ;
        RECT 1495.730 2941.090 1496.910 2942.270 ;
        RECT 1494.130 2939.490 1495.310 2940.670 ;
        RECT 1495.730 2939.490 1496.910 2940.670 ;
        RECT 1494.130 2761.090 1495.310 2762.270 ;
        RECT 1495.730 2761.090 1496.910 2762.270 ;
        RECT 1494.130 2759.490 1495.310 2760.670 ;
        RECT 1495.730 2759.490 1496.910 2760.670 ;
        RECT 1494.130 2581.090 1495.310 2582.270 ;
        RECT 1495.730 2581.090 1496.910 2582.270 ;
        RECT 1494.130 2579.490 1495.310 2580.670 ;
        RECT 1495.730 2579.490 1496.910 2580.670 ;
        RECT 1494.130 2401.090 1495.310 2402.270 ;
        RECT 1495.730 2401.090 1496.910 2402.270 ;
        RECT 1494.130 2399.490 1495.310 2400.670 ;
        RECT 1495.730 2399.490 1496.910 2400.670 ;
        RECT 1494.130 2221.090 1495.310 2222.270 ;
        RECT 1495.730 2221.090 1496.910 2222.270 ;
        RECT 1494.130 2219.490 1495.310 2220.670 ;
        RECT 1495.730 2219.490 1496.910 2220.670 ;
        RECT 1494.130 2041.090 1495.310 2042.270 ;
        RECT 1495.730 2041.090 1496.910 2042.270 ;
        RECT 1494.130 2039.490 1495.310 2040.670 ;
        RECT 1495.730 2039.490 1496.910 2040.670 ;
        RECT 1494.130 1861.090 1495.310 1862.270 ;
        RECT 1495.730 1861.090 1496.910 1862.270 ;
        RECT 1494.130 1859.490 1495.310 1860.670 ;
        RECT 1495.730 1859.490 1496.910 1860.670 ;
        RECT 1494.130 1681.090 1495.310 1682.270 ;
        RECT 1495.730 1681.090 1496.910 1682.270 ;
        RECT 1494.130 1679.490 1495.310 1680.670 ;
        RECT 1495.730 1679.490 1496.910 1680.670 ;
        RECT 1494.130 1501.090 1495.310 1502.270 ;
        RECT 1495.730 1501.090 1496.910 1502.270 ;
        RECT 1494.130 1499.490 1495.310 1500.670 ;
        RECT 1495.730 1499.490 1496.910 1500.670 ;
        RECT 1494.130 1321.090 1495.310 1322.270 ;
        RECT 1495.730 1321.090 1496.910 1322.270 ;
        RECT 1494.130 1319.490 1495.310 1320.670 ;
        RECT 1495.730 1319.490 1496.910 1320.670 ;
        RECT 1494.130 1141.090 1495.310 1142.270 ;
        RECT 1495.730 1141.090 1496.910 1142.270 ;
        RECT 1494.130 1139.490 1495.310 1140.670 ;
        RECT 1495.730 1139.490 1496.910 1140.670 ;
        RECT 1494.130 961.090 1495.310 962.270 ;
        RECT 1495.730 961.090 1496.910 962.270 ;
        RECT 1494.130 959.490 1495.310 960.670 ;
        RECT 1495.730 959.490 1496.910 960.670 ;
        RECT 1494.130 781.090 1495.310 782.270 ;
        RECT 1495.730 781.090 1496.910 782.270 ;
        RECT 1494.130 779.490 1495.310 780.670 ;
        RECT 1495.730 779.490 1496.910 780.670 ;
        RECT 1494.130 601.090 1495.310 602.270 ;
        RECT 1495.730 601.090 1496.910 602.270 ;
        RECT 1494.130 599.490 1495.310 600.670 ;
        RECT 1495.730 599.490 1496.910 600.670 ;
        RECT 1494.130 421.090 1495.310 422.270 ;
        RECT 1495.730 421.090 1496.910 422.270 ;
        RECT 1494.130 419.490 1495.310 420.670 ;
        RECT 1495.730 419.490 1496.910 420.670 ;
        RECT 1494.130 241.090 1495.310 242.270 ;
        RECT 1495.730 241.090 1496.910 242.270 ;
        RECT 1494.130 239.490 1495.310 240.670 ;
        RECT 1495.730 239.490 1496.910 240.670 ;
        RECT 1494.130 61.090 1495.310 62.270 ;
        RECT 1495.730 61.090 1496.910 62.270 ;
        RECT 1494.130 59.490 1495.310 60.670 ;
        RECT 1495.730 59.490 1496.910 60.670 ;
        RECT 1494.130 -14.060 1495.310 -12.880 ;
        RECT 1495.730 -14.060 1496.910 -12.880 ;
        RECT 1494.130 -15.660 1495.310 -14.480 ;
        RECT 1495.730 -15.660 1496.910 -14.480 ;
        RECT 1674.130 3534.160 1675.310 3535.340 ;
        RECT 1675.730 3534.160 1676.910 3535.340 ;
        RECT 1674.130 3532.560 1675.310 3533.740 ;
        RECT 1675.730 3532.560 1676.910 3533.740 ;
        RECT 1674.130 3481.090 1675.310 3482.270 ;
        RECT 1675.730 3481.090 1676.910 3482.270 ;
        RECT 1674.130 3479.490 1675.310 3480.670 ;
        RECT 1675.730 3479.490 1676.910 3480.670 ;
        RECT 1674.130 3301.090 1675.310 3302.270 ;
        RECT 1675.730 3301.090 1676.910 3302.270 ;
        RECT 1674.130 3299.490 1675.310 3300.670 ;
        RECT 1675.730 3299.490 1676.910 3300.670 ;
        RECT 1674.130 3121.090 1675.310 3122.270 ;
        RECT 1675.730 3121.090 1676.910 3122.270 ;
        RECT 1674.130 3119.490 1675.310 3120.670 ;
        RECT 1675.730 3119.490 1676.910 3120.670 ;
        RECT 1674.130 2941.090 1675.310 2942.270 ;
        RECT 1675.730 2941.090 1676.910 2942.270 ;
        RECT 1674.130 2939.490 1675.310 2940.670 ;
        RECT 1675.730 2939.490 1676.910 2940.670 ;
        RECT 1674.130 2761.090 1675.310 2762.270 ;
        RECT 1675.730 2761.090 1676.910 2762.270 ;
        RECT 1674.130 2759.490 1675.310 2760.670 ;
        RECT 1675.730 2759.490 1676.910 2760.670 ;
        RECT 1674.130 2581.090 1675.310 2582.270 ;
        RECT 1675.730 2581.090 1676.910 2582.270 ;
        RECT 1674.130 2579.490 1675.310 2580.670 ;
        RECT 1675.730 2579.490 1676.910 2580.670 ;
        RECT 1674.130 2401.090 1675.310 2402.270 ;
        RECT 1675.730 2401.090 1676.910 2402.270 ;
        RECT 1674.130 2399.490 1675.310 2400.670 ;
        RECT 1675.730 2399.490 1676.910 2400.670 ;
        RECT 1674.130 2221.090 1675.310 2222.270 ;
        RECT 1675.730 2221.090 1676.910 2222.270 ;
        RECT 1674.130 2219.490 1675.310 2220.670 ;
        RECT 1675.730 2219.490 1676.910 2220.670 ;
        RECT 1674.130 2041.090 1675.310 2042.270 ;
        RECT 1675.730 2041.090 1676.910 2042.270 ;
        RECT 1674.130 2039.490 1675.310 2040.670 ;
        RECT 1675.730 2039.490 1676.910 2040.670 ;
        RECT 1674.130 1861.090 1675.310 1862.270 ;
        RECT 1675.730 1861.090 1676.910 1862.270 ;
        RECT 1674.130 1859.490 1675.310 1860.670 ;
        RECT 1675.730 1859.490 1676.910 1860.670 ;
        RECT 1674.130 1681.090 1675.310 1682.270 ;
        RECT 1675.730 1681.090 1676.910 1682.270 ;
        RECT 1674.130 1679.490 1675.310 1680.670 ;
        RECT 1675.730 1679.490 1676.910 1680.670 ;
        RECT 1674.130 1501.090 1675.310 1502.270 ;
        RECT 1675.730 1501.090 1676.910 1502.270 ;
        RECT 1674.130 1499.490 1675.310 1500.670 ;
        RECT 1675.730 1499.490 1676.910 1500.670 ;
        RECT 1674.130 1321.090 1675.310 1322.270 ;
        RECT 1675.730 1321.090 1676.910 1322.270 ;
        RECT 1674.130 1319.490 1675.310 1320.670 ;
        RECT 1675.730 1319.490 1676.910 1320.670 ;
        RECT 1674.130 1141.090 1675.310 1142.270 ;
        RECT 1675.730 1141.090 1676.910 1142.270 ;
        RECT 1674.130 1139.490 1675.310 1140.670 ;
        RECT 1675.730 1139.490 1676.910 1140.670 ;
        RECT 1674.130 961.090 1675.310 962.270 ;
        RECT 1675.730 961.090 1676.910 962.270 ;
        RECT 1674.130 959.490 1675.310 960.670 ;
        RECT 1675.730 959.490 1676.910 960.670 ;
        RECT 1674.130 781.090 1675.310 782.270 ;
        RECT 1675.730 781.090 1676.910 782.270 ;
        RECT 1674.130 779.490 1675.310 780.670 ;
        RECT 1675.730 779.490 1676.910 780.670 ;
        RECT 1674.130 601.090 1675.310 602.270 ;
        RECT 1675.730 601.090 1676.910 602.270 ;
        RECT 1674.130 599.490 1675.310 600.670 ;
        RECT 1675.730 599.490 1676.910 600.670 ;
        RECT 1674.130 421.090 1675.310 422.270 ;
        RECT 1675.730 421.090 1676.910 422.270 ;
        RECT 1674.130 419.490 1675.310 420.670 ;
        RECT 1675.730 419.490 1676.910 420.670 ;
        RECT 1674.130 241.090 1675.310 242.270 ;
        RECT 1675.730 241.090 1676.910 242.270 ;
        RECT 1674.130 239.490 1675.310 240.670 ;
        RECT 1675.730 239.490 1676.910 240.670 ;
        RECT 1674.130 61.090 1675.310 62.270 ;
        RECT 1675.730 61.090 1676.910 62.270 ;
        RECT 1674.130 59.490 1675.310 60.670 ;
        RECT 1675.730 59.490 1676.910 60.670 ;
        RECT 1674.130 -14.060 1675.310 -12.880 ;
        RECT 1675.730 -14.060 1676.910 -12.880 ;
        RECT 1674.130 -15.660 1675.310 -14.480 ;
        RECT 1675.730 -15.660 1676.910 -14.480 ;
        RECT 1854.130 3534.160 1855.310 3535.340 ;
        RECT 1855.730 3534.160 1856.910 3535.340 ;
        RECT 1854.130 3532.560 1855.310 3533.740 ;
        RECT 1855.730 3532.560 1856.910 3533.740 ;
        RECT 1854.130 3481.090 1855.310 3482.270 ;
        RECT 1855.730 3481.090 1856.910 3482.270 ;
        RECT 1854.130 3479.490 1855.310 3480.670 ;
        RECT 1855.730 3479.490 1856.910 3480.670 ;
        RECT 1854.130 3301.090 1855.310 3302.270 ;
        RECT 1855.730 3301.090 1856.910 3302.270 ;
        RECT 1854.130 3299.490 1855.310 3300.670 ;
        RECT 1855.730 3299.490 1856.910 3300.670 ;
        RECT 1854.130 3121.090 1855.310 3122.270 ;
        RECT 1855.730 3121.090 1856.910 3122.270 ;
        RECT 1854.130 3119.490 1855.310 3120.670 ;
        RECT 1855.730 3119.490 1856.910 3120.670 ;
        RECT 1854.130 2941.090 1855.310 2942.270 ;
        RECT 1855.730 2941.090 1856.910 2942.270 ;
        RECT 1854.130 2939.490 1855.310 2940.670 ;
        RECT 1855.730 2939.490 1856.910 2940.670 ;
        RECT 1854.130 2761.090 1855.310 2762.270 ;
        RECT 1855.730 2761.090 1856.910 2762.270 ;
        RECT 1854.130 2759.490 1855.310 2760.670 ;
        RECT 1855.730 2759.490 1856.910 2760.670 ;
        RECT 1854.130 2581.090 1855.310 2582.270 ;
        RECT 1855.730 2581.090 1856.910 2582.270 ;
        RECT 1854.130 2579.490 1855.310 2580.670 ;
        RECT 1855.730 2579.490 1856.910 2580.670 ;
        RECT 1854.130 2401.090 1855.310 2402.270 ;
        RECT 1855.730 2401.090 1856.910 2402.270 ;
        RECT 1854.130 2399.490 1855.310 2400.670 ;
        RECT 1855.730 2399.490 1856.910 2400.670 ;
        RECT 1854.130 2221.090 1855.310 2222.270 ;
        RECT 1855.730 2221.090 1856.910 2222.270 ;
        RECT 1854.130 2219.490 1855.310 2220.670 ;
        RECT 1855.730 2219.490 1856.910 2220.670 ;
        RECT 1854.130 2041.090 1855.310 2042.270 ;
        RECT 1855.730 2041.090 1856.910 2042.270 ;
        RECT 1854.130 2039.490 1855.310 2040.670 ;
        RECT 1855.730 2039.490 1856.910 2040.670 ;
        RECT 1854.130 1861.090 1855.310 1862.270 ;
        RECT 1855.730 1861.090 1856.910 1862.270 ;
        RECT 1854.130 1859.490 1855.310 1860.670 ;
        RECT 1855.730 1859.490 1856.910 1860.670 ;
        RECT 1854.130 1681.090 1855.310 1682.270 ;
        RECT 1855.730 1681.090 1856.910 1682.270 ;
        RECT 1854.130 1679.490 1855.310 1680.670 ;
        RECT 1855.730 1679.490 1856.910 1680.670 ;
        RECT 1854.130 1501.090 1855.310 1502.270 ;
        RECT 1855.730 1501.090 1856.910 1502.270 ;
        RECT 1854.130 1499.490 1855.310 1500.670 ;
        RECT 1855.730 1499.490 1856.910 1500.670 ;
        RECT 1854.130 1321.090 1855.310 1322.270 ;
        RECT 1855.730 1321.090 1856.910 1322.270 ;
        RECT 1854.130 1319.490 1855.310 1320.670 ;
        RECT 1855.730 1319.490 1856.910 1320.670 ;
        RECT 1854.130 1141.090 1855.310 1142.270 ;
        RECT 1855.730 1141.090 1856.910 1142.270 ;
        RECT 1854.130 1139.490 1855.310 1140.670 ;
        RECT 1855.730 1139.490 1856.910 1140.670 ;
        RECT 1854.130 961.090 1855.310 962.270 ;
        RECT 1855.730 961.090 1856.910 962.270 ;
        RECT 1854.130 959.490 1855.310 960.670 ;
        RECT 1855.730 959.490 1856.910 960.670 ;
        RECT 1854.130 781.090 1855.310 782.270 ;
        RECT 1855.730 781.090 1856.910 782.270 ;
        RECT 1854.130 779.490 1855.310 780.670 ;
        RECT 1855.730 779.490 1856.910 780.670 ;
        RECT 1854.130 601.090 1855.310 602.270 ;
        RECT 1855.730 601.090 1856.910 602.270 ;
        RECT 1854.130 599.490 1855.310 600.670 ;
        RECT 1855.730 599.490 1856.910 600.670 ;
        RECT 1854.130 421.090 1855.310 422.270 ;
        RECT 1855.730 421.090 1856.910 422.270 ;
        RECT 1854.130 419.490 1855.310 420.670 ;
        RECT 1855.730 419.490 1856.910 420.670 ;
        RECT 1854.130 241.090 1855.310 242.270 ;
        RECT 1855.730 241.090 1856.910 242.270 ;
        RECT 1854.130 239.490 1855.310 240.670 ;
        RECT 1855.730 239.490 1856.910 240.670 ;
        RECT 1854.130 61.090 1855.310 62.270 ;
        RECT 1855.730 61.090 1856.910 62.270 ;
        RECT 1854.130 59.490 1855.310 60.670 ;
        RECT 1855.730 59.490 1856.910 60.670 ;
        RECT 1854.130 -14.060 1855.310 -12.880 ;
        RECT 1855.730 -14.060 1856.910 -12.880 ;
        RECT 1854.130 -15.660 1855.310 -14.480 ;
        RECT 1855.730 -15.660 1856.910 -14.480 ;
        RECT 2034.130 3534.160 2035.310 3535.340 ;
        RECT 2035.730 3534.160 2036.910 3535.340 ;
        RECT 2034.130 3532.560 2035.310 3533.740 ;
        RECT 2035.730 3532.560 2036.910 3533.740 ;
        RECT 2034.130 3481.090 2035.310 3482.270 ;
        RECT 2035.730 3481.090 2036.910 3482.270 ;
        RECT 2034.130 3479.490 2035.310 3480.670 ;
        RECT 2035.730 3479.490 2036.910 3480.670 ;
        RECT 2034.130 3301.090 2035.310 3302.270 ;
        RECT 2035.730 3301.090 2036.910 3302.270 ;
        RECT 2034.130 3299.490 2035.310 3300.670 ;
        RECT 2035.730 3299.490 2036.910 3300.670 ;
        RECT 2034.130 3121.090 2035.310 3122.270 ;
        RECT 2035.730 3121.090 2036.910 3122.270 ;
        RECT 2034.130 3119.490 2035.310 3120.670 ;
        RECT 2035.730 3119.490 2036.910 3120.670 ;
        RECT 2034.130 2941.090 2035.310 2942.270 ;
        RECT 2035.730 2941.090 2036.910 2942.270 ;
        RECT 2034.130 2939.490 2035.310 2940.670 ;
        RECT 2035.730 2939.490 2036.910 2940.670 ;
        RECT 2034.130 2761.090 2035.310 2762.270 ;
        RECT 2035.730 2761.090 2036.910 2762.270 ;
        RECT 2034.130 2759.490 2035.310 2760.670 ;
        RECT 2035.730 2759.490 2036.910 2760.670 ;
        RECT 2034.130 2581.090 2035.310 2582.270 ;
        RECT 2035.730 2581.090 2036.910 2582.270 ;
        RECT 2034.130 2579.490 2035.310 2580.670 ;
        RECT 2035.730 2579.490 2036.910 2580.670 ;
        RECT 2034.130 2401.090 2035.310 2402.270 ;
        RECT 2035.730 2401.090 2036.910 2402.270 ;
        RECT 2034.130 2399.490 2035.310 2400.670 ;
        RECT 2035.730 2399.490 2036.910 2400.670 ;
        RECT 2034.130 2221.090 2035.310 2222.270 ;
        RECT 2035.730 2221.090 2036.910 2222.270 ;
        RECT 2034.130 2219.490 2035.310 2220.670 ;
        RECT 2035.730 2219.490 2036.910 2220.670 ;
        RECT 2034.130 2041.090 2035.310 2042.270 ;
        RECT 2035.730 2041.090 2036.910 2042.270 ;
        RECT 2034.130 2039.490 2035.310 2040.670 ;
        RECT 2035.730 2039.490 2036.910 2040.670 ;
        RECT 2034.130 1861.090 2035.310 1862.270 ;
        RECT 2035.730 1861.090 2036.910 1862.270 ;
        RECT 2034.130 1859.490 2035.310 1860.670 ;
        RECT 2035.730 1859.490 2036.910 1860.670 ;
        RECT 2034.130 1681.090 2035.310 1682.270 ;
        RECT 2035.730 1681.090 2036.910 1682.270 ;
        RECT 2034.130 1679.490 2035.310 1680.670 ;
        RECT 2035.730 1679.490 2036.910 1680.670 ;
        RECT 2034.130 1501.090 2035.310 1502.270 ;
        RECT 2035.730 1501.090 2036.910 1502.270 ;
        RECT 2034.130 1499.490 2035.310 1500.670 ;
        RECT 2035.730 1499.490 2036.910 1500.670 ;
        RECT 2034.130 1321.090 2035.310 1322.270 ;
        RECT 2035.730 1321.090 2036.910 1322.270 ;
        RECT 2034.130 1319.490 2035.310 1320.670 ;
        RECT 2035.730 1319.490 2036.910 1320.670 ;
        RECT 2034.130 1141.090 2035.310 1142.270 ;
        RECT 2035.730 1141.090 2036.910 1142.270 ;
        RECT 2034.130 1139.490 2035.310 1140.670 ;
        RECT 2035.730 1139.490 2036.910 1140.670 ;
        RECT 2034.130 961.090 2035.310 962.270 ;
        RECT 2035.730 961.090 2036.910 962.270 ;
        RECT 2034.130 959.490 2035.310 960.670 ;
        RECT 2035.730 959.490 2036.910 960.670 ;
        RECT 2034.130 781.090 2035.310 782.270 ;
        RECT 2035.730 781.090 2036.910 782.270 ;
        RECT 2034.130 779.490 2035.310 780.670 ;
        RECT 2035.730 779.490 2036.910 780.670 ;
        RECT 2034.130 601.090 2035.310 602.270 ;
        RECT 2035.730 601.090 2036.910 602.270 ;
        RECT 2034.130 599.490 2035.310 600.670 ;
        RECT 2035.730 599.490 2036.910 600.670 ;
        RECT 2034.130 421.090 2035.310 422.270 ;
        RECT 2035.730 421.090 2036.910 422.270 ;
        RECT 2034.130 419.490 2035.310 420.670 ;
        RECT 2035.730 419.490 2036.910 420.670 ;
        RECT 2034.130 241.090 2035.310 242.270 ;
        RECT 2035.730 241.090 2036.910 242.270 ;
        RECT 2034.130 239.490 2035.310 240.670 ;
        RECT 2035.730 239.490 2036.910 240.670 ;
        RECT 2034.130 61.090 2035.310 62.270 ;
        RECT 2035.730 61.090 2036.910 62.270 ;
        RECT 2034.130 59.490 2035.310 60.670 ;
        RECT 2035.730 59.490 2036.910 60.670 ;
        RECT 2034.130 -14.060 2035.310 -12.880 ;
        RECT 2035.730 -14.060 2036.910 -12.880 ;
        RECT 2034.130 -15.660 2035.310 -14.480 ;
        RECT 2035.730 -15.660 2036.910 -14.480 ;
        RECT 2214.130 3534.160 2215.310 3535.340 ;
        RECT 2215.730 3534.160 2216.910 3535.340 ;
        RECT 2214.130 3532.560 2215.310 3533.740 ;
        RECT 2215.730 3532.560 2216.910 3533.740 ;
        RECT 2214.130 3481.090 2215.310 3482.270 ;
        RECT 2215.730 3481.090 2216.910 3482.270 ;
        RECT 2214.130 3479.490 2215.310 3480.670 ;
        RECT 2215.730 3479.490 2216.910 3480.670 ;
        RECT 2214.130 3301.090 2215.310 3302.270 ;
        RECT 2215.730 3301.090 2216.910 3302.270 ;
        RECT 2214.130 3299.490 2215.310 3300.670 ;
        RECT 2215.730 3299.490 2216.910 3300.670 ;
        RECT 2214.130 3121.090 2215.310 3122.270 ;
        RECT 2215.730 3121.090 2216.910 3122.270 ;
        RECT 2214.130 3119.490 2215.310 3120.670 ;
        RECT 2215.730 3119.490 2216.910 3120.670 ;
        RECT 2214.130 2941.090 2215.310 2942.270 ;
        RECT 2215.730 2941.090 2216.910 2942.270 ;
        RECT 2214.130 2939.490 2215.310 2940.670 ;
        RECT 2215.730 2939.490 2216.910 2940.670 ;
        RECT 2214.130 2761.090 2215.310 2762.270 ;
        RECT 2215.730 2761.090 2216.910 2762.270 ;
        RECT 2214.130 2759.490 2215.310 2760.670 ;
        RECT 2215.730 2759.490 2216.910 2760.670 ;
        RECT 2214.130 2581.090 2215.310 2582.270 ;
        RECT 2215.730 2581.090 2216.910 2582.270 ;
        RECT 2214.130 2579.490 2215.310 2580.670 ;
        RECT 2215.730 2579.490 2216.910 2580.670 ;
        RECT 2214.130 2401.090 2215.310 2402.270 ;
        RECT 2215.730 2401.090 2216.910 2402.270 ;
        RECT 2214.130 2399.490 2215.310 2400.670 ;
        RECT 2215.730 2399.490 2216.910 2400.670 ;
        RECT 2214.130 2221.090 2215.310 2222.270 ;
        RECT 2215.730 2221.090 2216.910 2222.270 ;
        RECT 2214.130 2219.490 2215.310 2220.670 ;
        RECT 2215.730 2219.490 2216.910 2220.670 ;
        RECT 2214.130 2041.090 2215.310 2042.270 ;
        RECT 2215.730 2041.090 2216.910 2042.270 ;
        RECT 2214.130 2039.490 2215.310 2040.670 ;
        RECT 2215.730 2039.490 2216.910 2040.670 ;
        RECT 2214.130 1861.090 2215.310 1862.270 ;
        RECT 2215.730 1861.090 2216.910 1862.270 ;
        RECT 2214.130 1859.490 2215.310 1860.670 ;
        RECT 2215.730 1859.490 2216.910 1860.670 ;
        RECT 2214.130 1681.090 2215.310 1682.270 ;
        RECT 2215.730 1681.090 2216.910 1682.270 ;
        RECT 2214.130 1679.490 2215.310 1680.670 ;
        RECT 2215.730 1679.490 2216.910 1680.670 ;
        RECT 2214.130 1501.090 2215.310 1502.270 ;
        RECT 2215.730 1501.090 2216.910 1502.270 ;
        RECT 2214.130 1499.490 2215.310 1500.670 ;
        RECT 2215.730 1499.490 2216.910 1500.670 ;
        RECT 2214.130 1321.090 2215.310 1322.270 ;
        RECT 2215.730 1321.090 2216.910 1322.270 ;
        RECT 2214.130 1319.490 2215.310 1320.670 ;
        RECT 2215.730 1319.490 2216.910 1320.670 ;
        RECT 2214.130 1141.090 2215.310 1142.270 ;
        RECT 2215.730 1141.090 2216.910 1142.270 ;
        RECT 2214.130 1139.490 2215.310 1140.670 ;
        RECT 2215.730 1139.490 2216.910 1140.670 ;
        RECT 2214.130 961.090 2215.310 962.270 ;
        RECT 2215.730 961.090 2216.910 962.270 ;
        RECT 2214.130 959.490 2215.310 960.670 ;
        RECT 2215.730 959.490 2216.910 960.670 ;
        RECT 2214.130 781.090 2215.310 782.270 ;
        RECT 2215.730 781.090 2216.910 782.270 ;
        RECT 2214.130 779.490 2215.310 780.670 ;
        RECT 2215.730 779.490 2216.910 780.670 ;
        RECT 2214.130 601.090 2215.310 602.270 ;
        RECT 2215.730 601.090 2216.910 602.270 ;
        RECT 2214.130 599.490 2215.310 600.670 ;
        RECT 2215.730 599.490 2216.910 600.670 ;
        RECT 2214.130 421.090 2215.310 422.270 ;
        RECT 2215.730 421.090 2216.910 422.270 ;
        RECT 2214.130 419.490 2215.310 420.670 ;
        RECT 2215.730 419.490 2216.910 420.670 ;
        RECT 2214.130 241.090 2215.310 242.270 ;
        RECT 2215.730 241.090 2216.910 242.270 ;
        RECT 2214.130 239.490 2215.310 240.670 ;
        RECT 2215.730 239.490 2216.910 240.670 ;
        RECT 2214.130 61.090 2215.310 62.270 ;
        RECT 2215.730 61.090 2216.910 62.270 ;
        RECT 2214.130 59.490 2215.310 60.670 ;
        RECT 2215.730 59.490 2216.910 60.670 ;
        RECT 2214.130 -14.060 2215.310 -12.880 ;
        RECT 2215.730 -14.060 2216.910 -12.880 ;
        RECT 2214.130 -15.660 2215.310 -14.480 ;
        RECT 2215.730 -15.660 2216.910 -14.480 ;
        RECT 2394.130 3534.160 2395.310 3535.340 ;
        RECT 2395.730 3534.160 2396.910 3535.340 ;
        RECT 2394.130 3532.560 2395.310 3533.740 ;
        RECT 2395.730 3532.560 2396.910 3533.740 ;
        RECT 2394.130 3481.090 2395.310 3482.270 ;
        RECT 2395.730 3481.090 2396.910 3482.270 ;
        RECT 2394.130 3479.490 2395.310 3480.670 ;
        RECT 2395.730 3479.490 2396.910 3480.670 ;
        RECT 2394.130 3301.090 2395.310 3302.270 ;
        RECT 2395.730 3301.090 2396.910 3302.270 ;
        RECT 2394.130 3299.490 2395.310 3300.670 ;
        RECT 2395.730 3299.490 2396.910 3300.670 ;
        RECT 2394.130 3121.090 2395.310 3122.270 ;
        RECT 2395.730 3121.090 2396.910 3122.270 ;
        RECT 2394.130 3119.490 2395.310 3120.670 ;
        RECT 2395.730 3119.490 2396.910 3120.670 ;
        RECT 2394.130 2941.090 2395.310 2942.270 ;
        RECT 2395.730 2941.090 2396.910 2942.270 ;
        RECT 2394.130 2939.490 2395.310 2940.670 ;
        RECT 2395.730 2939.490 2396.910 2940.670 ;
        RECT 2394.130 2761.090 2395.310 2762.270 ;
        RECT 2395.730 2761.090 2396.910 2762.270 ;
        RECT 2394.130 2759.490 2395.310 2760.670 ;
        RECT 2395.730 2759.490 2396.910 2760.670 ;
        RECT 2394.130 2581.090 2395.310 2582.270 ;
        RECT 2395.730 2581.090 2396.910 2582.270 ;
        RECT 2394.130 2579.490 2395.310 2580.670 ;
        RECT 2395.730 2579.490 2396.910 2580.670 ;
        RECT 2394.130 2401.090 2395.310 2402.270 ;
        RECT 2395.730 2401.090 2396.910 2402.270 ;
        RECT 2394.130 2399.490 2395.310 2400.670 ;
        RECT 2395.730 2399.490 2396.910 2400.670 ;
        RECT 2394.130 2221.090 2395.310 2222.270 ;
        RECT 2395.730 2221.090 2396.910 2222.270 ;
        RECT 2394.130 2219.490 2395.310 2220.670 ;
        RECT 2395.730 2219.490 2396.910 2220.670 ;
        RECT 2394.130 2041.090 2395.310 2042.270 ;
        RECT 2395.730 2041.090 2396.910 2042.270 ;
        RECT 2394.130 2039.490 2395.310 2040.670 ;
        RECT 2395.730 2039.490 2396.910 2040.670 ;
        RECT 2394.130 1861.090 2395.310 1862.270 ;
        RECT 2395.730 1861.090 2396.910 1862.270 ;
        RECT 2394.130 1859.490 2395.310 1860.670 ;
        RECT 2395.730 1859.490 2396.910 1860.670 ;
        RECT 2394.130 1681.090 2395.310 1682.270 ;
        RECT 2395.730 1681.090 2396.910 1682.270 ;
        RECT 2394.130 1679.490 2395.310 1680.670 ;
        RECT 2395.730 1679.490 2396.910 1680.670 ;
        RECT 2394.130 1501.090 2395.310 1502.270 ;
        RECT 2395.730 1501.090 2396.910 1502.270 ;
        RECT 2394.130 1499.490 2395.310 1500.670 ;
        RECT 2395.730 1499.490 2396.910 1500.670 ;
        RECT 2394.130 1321.090 2395.310 1322.270 ;
        RECT 2395.730 1321.090 2396.910 1322.270 ;
        RECT 2394.130 1319.490 2395.310 1320.670 ;
        RECT 2395.730 1319.490 2396.910 1320.670 ;
        RECT 2394.130 1141.090 2395.310 1142.270 ;
        RECT 2395.730 1141.090 2396.910 1142.270 ;
        RECT 2394.130 1139.490 2395.310 1140.670 ;
        RECT 2395.730 1139.490 2396.910 1140.670 ;
        RECT 2394.130 961.090 2395.310 962.270 ;
        RECT 2395.730 961.090 2396.910 962.270 ;
        RECT 2394.130 959.490 2395.310 960.670 ;
        RECT 2395.730 959.490 2396.910 960.670 ;
        RECT 2394.130 781.090 2395.310 782.270 ;
        RECT 2395.730 781.090 2396.910 782.270 ;
        RECT 2394.130 779.490 2395.310 780.670 ;
        RECT 2395.730 779.490 2396.910 780.670 ;
        RECT 2394.130 601.090 2395.310 602.270 ;
        RECT 2395.730 601.090 2396.910 602.270 ;
        RECT 2394.130 599.490 2395.310 600.670 ;
        RECT 2395.730 599.490 2396.910 600.670 ;
        RECT 2394.130 421.090 2395.310 422.270 ;
        RECT 2395.730 421.090 2396.910 422.270 ;
        RECT 2394.130 419.490 2395.310 420.670 ;
        RECT 2395.730 419.490 2396.910 420.670 ;
        RECT 2394.130 241.090 2395.310 242.270 ;
        RECT 2395.730 241.090 2396.910 242.270 ;
        RECT 2394.130 239.490 2395.310 240.670 ;
        RECT 2395.730 239.490 2396.910 240.670 ;
        RECT 2394.130 61.090 2395.310 62.270 ;
        RECT 2395.730 61.090 2396.910 62.270 ;
        RECT 2394.130 59.490 2395.310 60.670 ;
        RECT 2395.730 59.490 2396.910 60.670 ;
        RECT 2394.130 -14.060 2395.310 -12.880 ;
        RECT 2395.730 -14.060 2396.910 -12.880 ;
        RECT 2394.130 -15.660 2395.310 -14.480 ;
        RECT 2395.730 -15.660 2396.910 -14.480 ;
        RECT 2574.130 3534.160 2575.310 3535.340 ;
        RECT 2575.730 3534.160 2576.910 3535.340 ;
        RECT 2574.130 3532.560 2575.310 3533.740 ;
        RECT 2575.730 3532.560 2576.910 3533.740 ;
        RECT 2574.130 3481.090 2575.310 3482.270 ;
        RECT 2575.730 3481.090 2576.910 3482.270 ;
        RECT 2574.130 3479.490 2575.310 3480.670 ;
        RECT 2575.730 3479.490 2576.910 3480.670 ;
        RECT 2574.130 3301.090 2575.310 3302.270 ;
        RECT 2575.730 3301.090 2576.910 3302.270 ;
        RECT 2574.130 3299.490 2575.310 3300.670 ;
        RECT 2575.730 3299.490 2576.910 3300.670 ;
        RECT 2574.130 3121.090 2575.310 3122.270 ;
        RECT 2575.730 3121.090 2576.910 3122.270 ;
        RECT 2574.130 3119.490 2575.310 3120.670 ;
        RECT 2575.730 3119.490 2576.910 3120.670 ;
        RECT 2574.130 2941.090 2575.310 2942.270 ;
        RECT 2575.730 2941.090 2576.910 2942.270 ;
        RECT 2574.130 2939.490 2575.310 2940.670 ;
        RECT 2575.730 2939.490 2576.910 2940.670 ;
        RECT 2574.130 2761.090 2575.310 2762.270 ;
        RECT 2575.730 2761.090 2576.910 2762.270 ;
        RECT 2574.130 2759.490 2575.310 2760.670 ;
        RECT 2575.730 2759.490 2576.910 2760.670 ;
        RECT 2574.130 2581.090 2575.310 2582.270 ;
        RECT 2575.730 2581.090 2576.910 2582.270 ;
        RECT 2574.130 2579.490 2575.310 2580.670 ;
        RECT 2575.730 2579.490 2576.910 2580.670 ;
        RECT 2574.130 2401.090 2575.310 2402.270 ;
        RECT 2575.730 2401.090 2576.910 2402.270 ;
        RECT 2574.130 2399.490 2575.310 2400.670 ;
        RECT 2575.730 2399.490 2576.910 2400.670 ;
        RECT 2574.130 2221.090 2575.310 2222.270 ;
        RECT 2575.730 2221.090 2576.910 2222.270 ;
        RECT 2574.130 2219.490 2575.310 2220.670 ;
        RECT 2575.730 2219.490 2576.910 2220.670 ;
        RECT 2574.130 2041.090 2575.310 2042.270 ;
        RECT 2575.730 2041.090 2576.910 2042.270 ;
        RECT 2574.130 2039.490 2575.310 2040.670 ;
        RECT 2575.730 2039.490 2576.910 2040.670 ;
        RECT 2574.130 1861.090 2575.310 1862.270 ;
        RECT 2575.730 1861.090 2576.910 1862.270 ;
        RECT 2574.130 1859.490 2575.310 1860.670 ;
        RECT 2575.730 1859.490 2576.910 1860.670 ;
        RECT 2574.130 1681.090 2575.310 1682.270 ;
        RECT 2575.730 1681.090 2576.910 1682.270 ;
        RECT 2574.130 1679.490 2575.310 1680.670 ;
        RECT 2575.730 1679.490 2576.910 1680.670 ;
        RECT 2574.130 1501.090 2575.310 1502.270 ;
        RECT 2575.730 1501.090 2576.910 1502.270 ;
        RECT 2574.130 1499.490 2575.310 1500.670 ;
        RECT 2575.730 1499.490 2576.910 1500.670 ;
        RECT 2574.130 1321.090 2575.310 1322.270 ;
        RECT 2575.730 1321.090 2576.910 1322.270 ;
        RECT 2574.130 1319.490 2575.310 1320.670 ;
        RECT 2575.730 1319.490 2576.910 1320.670 ;
        RECT 2574.130 1141.090 2575.310 1142.270 ;
        RECT 2575.730 1141.090 2576.910 1142.270 ;
        RECT 2574.130 1139.490 2575.310 1140.670 ;
        RECT 2575.730 1139.490 2576.910 1140.670 ;
        RECT 2574.130 961.090 2575.310 962.270 ;
        RECT 2575.730 961.090 2576.910 962.270 ;
        RECT 2574.130 959.490 2575.310 960.670 ;
        RECT 2575.730 959.490 2576.910 960.670 ;
        RECT 2574.130 781.090 2575.310 782.270 ;
        RECT 2575.730 781.090 2576.910 782.270 ;
        RECT 2574.130 779.490 2575.310 780.670 ;
        RECT 2575.730 779.490 2576.910 780.670 ;
        RECT 2574.130 601.090 2575.310 602.270 ;
        RECT 2575.730 601.090 2576.910 602.270 ;
        RECT 2574.130 599.490 2575.310 600.670 ;
        RECT 2575.730 599.490 2576.910 600.670 ;
        RECT 2574.130 421.090 2575.310 422.270 ;
        RECT 2575.730 421.090 2576.910 422.270 ;
        RECT 2574.130 419.490 2575.310 420.670 ;
        RECT 2575.730 419.490 2576.910 420.670 ;
        RECT 2574.130 241.090 2575.310 242.270 ;
        RECT 2575.730 241.090 2576.910 242.270 ;
        RECT 2574.130 239.490 2575.310 240.670 ;
        RECT 2575.730 239.490 2576.910 240.670 ;
        RECT 2574.130 61.090 2575.310 62.270 ;
        RECT 2575.730 61.090 2576.910 62.270 ;
        RECT 2574.130 59.490 2575.310 60.670 ;
        RECT 2575.730 59.490 2576.910 60.670 ;
        RECT 2574.130 -14.060 2575.310 -12.880 ;
        RECT 2575.730 -14.060 2576.910 -12.880 ;
        RECT 2574.130 -15.660 2575.310 -14.480 ;
        RECT 2575.730 -15.660 2576.910 -14.480 ;
        RECT 2754.130 3534.160 2755.310 3535.340 ;
        RECT 2755.730 3534.160 2756.910 3535.340 ;
        RECT 2754.130 3532.560 2755.310 3533.740 ;
        RECT 2755.730 3532.560 2756.910 3533.740 ;
        RECT 2754.130 3481.090 2755.310 3482.270 ;
        RECT 2755.730 3481.090 2756.910 3482.270 ;
        RECT 2754.130 3479.490 2755.310 3480.670 ;
        RECT 2755.730 3479.490 2756.910 3480.670 ;
        RECT 2754.130 3301.090 2755.310 3302.270 ;
        RECT 2755.730 3301.090 2756.910 3302.270 ;
        RECT 2754.130 3299.490 2755.310 3300.670 ;
        RECT 2755.730 3299.490 2756.910 3300.670 ;
        RECT 2754.130 3121.090 2755.310 3122.270 ;
        RECT 2755.730 3121.090 2756.910 3122.270 ;
        RECT 2754.130 3119.490 2755.310 3120.670 ;
        RECT 2755.730 3119.490 2756.910 3120.670 ;
        RECT 2754.130 2941.090 2755.310 2942.270 ;
        RECT 2755.730 2941.090 2756.910 2942.270 ;
        RECT 2754.130 2939.490 2755.310 2940.670 ;
        RECT 2755.730 2939.490 2756.910 2940.670 ;
        RECT 2754.130 2761.090 2755.310 2762.270 ;
        RECT 2755.730 2761.090 2756.910 2762.270 ;
        RECT 2754.130 2759.490 2755.310 2760.670 ;
        RECT 2755.730 2759.490 2756.910 2760.670 ;
        RECT 2754.130 2581.090 2755.310 2582.270 ;
        RECT 2755.730 2581.090 2756.910 2582.270 ;
        RECT 2754.130 2579.490 2755.310 2580.670 ;
        RECT 2755.730 2579.490 2756.910 2580.670 ;
        RECT 2754.130 2401.090 2755.310 2402.270 ;
        RECT 2755.730 2401.090 2756.910 2402.270 ;
        RECT 2754.130 2399.490 2755.310 2400.670 ;
        RECT 2755.730 2399.490 2756.910 2400.670 ;
        RECT 2754.130 2221.090 2755.310 2222.270 ;
        RECT 2755.730 2221.090 2756.910 2222.270 ;
        RECT 2754.130 2219.490 2755.310 2220.670 ;
        RECT 2755.730 2219.490 2756.910 2220.670 ;
        RECT 2754.130 2041.090 2755.310 2042.270 ;
        RECT 2755.730 2041.090 2756.910 2042.270 ;
        RECT 2754.130 2039.490 2755.310 2040.670 ;
        RECT 2755.730 2039.490 2756.910 2040.670 ;
        RECT 2754.130 1861.090 2755.310 1862.270 ;
        RECT 2755.730 1861.090 2756.910 1862.270 ;
        RECT 2754.130 1859.490 2755.310 1860.670 ;
        RECT 2755.730 1859.490 2756.910 1860.670 ;
        RECT 2754.130 1681.090 2755.310 1682.270 ;
        RECT 2755.730 1681.090 2756.910 1682.270 ;
        RECT 2754.130 1679.490 2755.310 1680.670 ;
        RECT 2755.730 1679.490 2756.910 1680.670 ;
        RECT 2754.130 1501.090 2755.310 1502.270 ;
        RECT 2755.730 1501.090 2756.910 1502.270 ;
        RECT 2754.130 1499.490 2755.310 1500.670 ;
        RECT 2755.730 1499.490 2756.910 1500.670 ;
        RECT 2754.130 1321.090 2755.310 1322.270 ;
        RECT 2755.730 1321.090 2756.910 1322.270 ;
        RECT 2754.130 1319.490 2755.310 1320.670 ;
        RECT 2755.730 1319.490 2756.910 1320.670 ;
        RECT 2754.130 1141.090 2755.310 1142.270 ;
        RECT 2755.730 1141.090 2756.910 1142.270 ;
        RECT 2754.130 1139.490 2755.310 1140.670 ;
        RECT 2755.730 1139.490 2756.910 1140.670 ;
        RECT 2754.130 961.090 2755.310 962.270 ;
        RECT 2755.730 961.090 2756.910 962.270 ;
        RECT 2754.130 959.490 2755.310 960.670 ;
        RECT 2755.730 959.490 2756.910 960.670 ;
        RECT 2754.130 781.090 2755.310 782.270 ;
        RECT 2755.730 781.090 2756.910 782.270 ;
        RECT 2754.130 779.490 2755.310 780.670 ;
        RECT 2755.730 779.490 2756.910 780.670 ;
        RECT 2754.130 601.090 2755.310 602.270 ;
        RECT 2755.730 601.090 2756.910 602.270 ;
        RECT 2754.130 599.490 2755.310 600.670 ;
        RECT 2755.730 599.490 2756.910 600.670 ;
        RECT 2754.130 421.090 2755.310 422.270 ;
        RECT 2755.730 421.090 2756.910 422.270 ;
        RECT 2754.130 419.490 2755.310 420.670 ;
        RECT 2755.730 419.490 2756.910 420.670 ;
        RECT 2754.130 241.090 2755.310 242.270 ;
        RECT 2755.730 241.090 2756.910 242.270 ;
        RECT 2754.130 239.490 2755.310 240.670 ;
        RECT 2755.730 239.490 2756.910 240.670 ;
        RECT 2754.130 61.090 2755.310 62.270 ;
        RECT 2755.730 61.090 2756.910 62.270 ;
        RECT 2754.130 59.490 2755.310 60.670 ;
        RECT 2755.730 59.490 2756.910 60.670 ;
        RECT 2754.130 -14.060 2755.310 -12.880 ;
        RECT 2755.730 -14.060 2756.910 -12.880 ;
        RECT 2754.130 -15.660 2755.310 -14.480 ;
        RECT 2755.730 -15.660 2756.910 -14.480 ;
        RECT 2937.860 3534.160 2939.040 3535.340 ;
        RECT 2939.460 3534.160 2940.640 3535.340 ;
        RECT 2937.860 3532.560 2939.040 3533.740 ;
        RECT 2939.460 3532.560 2940.640 3533.740 ;
        RECT 2937.860 3481.090 2939.040 3482.270 ;
        RECT 2939.460 3481.090 2940.640 3482.270 ;
        RECT 2937.860 3479.490 2939.040 3480.670 ;
        RECT 2939.460 3479.490 2940.640 3480.670 ;
        RECT 2937.860 3301.090 2939.040 3302.270 ;
        RECT 2939.460 3301.090 2940.640 3302.270 ;
        RECT 2937.860 3299.490 2939.040 3300.670 ;
        RECT 2939.460 3299.490 2940.640 3300.670 ;
        RECT 2937.860 3121.090 2939.040 3122.270 ;
        RECT 2939.460 3121.090 2940.640 3122.270 ;
        RECT 2937.860 3119.490 2939.040 3120.670 ;
        RECT 2939.460 3119.490 2940.640 3120.670 ;
        RECT 2937.860 2941.090 2939.040 2942.270 ;
        RECT 2939.460 2941.090 2940.640 2942.270 ;
        RECT 2937.860 2939.490 2939.040 2940.670 ;
        RECT 2939.460 2939.490 2940.640 2940.670 ;
        RECT 2937.860 2761.090 2939.040 2762.270 ;
        RECT 2939.460 2761.090 2940.640 2762.270 ;
        RECT 2937.860 2759.490 2939.040 2760.670 ;
        RECT 2939.460 2759.490 2940.640 2760.670 ;
        RECT 2937.860 2581.090 2939.040 2582.270 ;
        RECT 2939.460 2581.090 2940.640 2582.270 ;
        RECT 2937.860 2579.490 2939.040 2580.670 ;
        RECT 2939.460 2579.490 2940.640 2580.670 ;
        RECT 2937.860 2401.090 2939.040 2402.270 ;
        RECT 2939.460 2401.090 2940.640 2402.270 ;
        RECT 2937.860 2399.490 2939.040 2400.670 ;
        RECT 2939.460 2399.490 2940.640 2400.670 ;
        RECT 2937.860 2221.090 2939.040 2222.270 ;
        RECT 2939.460 2221.090 2940.640 2222.270 ;
        RECT 2937.860 2219.490 2939.040 2220.670 ;
        RECT 2939.460 2219.490 2940.640 2220.670 ;
        RECT 2937.860 2041.090 2939.040 2042.270 ;
        RECT 2939.460 2041.090 2940.640 2042.270 ;
        RECT 2937.860 2039.490 2939.040 2040.670 ;
        RECT 2939.460 2039.490 2940.640 2040.670 ;
        RECT 2937.860 1861.090 2939.040 1862.270 ;
        RECT 2939.460 1861.090 2940.640 1862.270 ;
        RECT 2937.860 1859.490 2939.040 1860.670 ;
        RECT 2939.460 1859.490 2940.640 1860.670 ;
        RECT 2937.860 1681.090 2939.040 1682.270 ;
        RECT 2939.460 1681.090 2940.640 1682.270 ;
        RECT 2937.860 1679.490 2939.040 1680.670 ;
        RECT 2939.460 1679.490 2940.640 1680.670 ;
        RECT 2937.860 1501.090 2939.040 1502.270 ;
        RECT 2939.460 1501.090 2940.640 1502.270 ;
        RECT 2937.860 1499.490 2939.040 1500.670 ;
        RECT 2939.460 1499.490 2940.640 1500.670 ;
        RECT 2937.860 1321.090 2939.040 1322.270 ;
        RECT 2939.460 1321.090 2940.640 1322.270 ;
        RECT 2937.860 1319.490 2939.040 1320.670 ;
        RECT 2939.460 1319.490 2940.640 1320.670 ;
        RECT 2937.860 1141.090 2939.040 1142.270 ;
        RECT 2939.460 1141.090 2940.640 1142.270 ;
        RECT 2937.860 1139.490 2939.040 1140.670 ;
        RECT 2939.460 1139.490 2940.640 1140.670 ;
        RECT 2937.860 961.090 2939.040 962.270 ;
        RECT 2939.460 961.090 2940.640 962.270 ;
        RECT 2937.860 959.490 2939.040 960.670 ;
        RECT 2939.460 959.490 2940.640 960.670 ;
        RECT 2937.860 781.090 2939.040 782.270 ;
        RECT 2939.460 781.090 2940.640 782.270 ;
        RECT 2937.860 779.490 2939.040 780.670 ;
        RECT 2939.460 779.490 2940.640 780.670 ;
        RECT 2937.860 601.090 2939.040 602.270 ;
        RECT 2939.460 601.090 2940.640 602.270 ;
        RECT 2937.860 599.490 2939.040 600.670 ;
        RECT 2939.460 599.490 2940.640 600.670 ;
        RECT 2937.860 421.090 2939.040 422.270 ;
        RECT 2939.460 421.090 2940.640 422.270 ;
        RECT 2937.860 419.490 2939.040 420.670 ;
        RECT 2939.460 419.490 2940.640 420.670 ;
        RECT 2937.860 241.090 2939.040 242.270 ;
        RECT 2939.460 241.090 2940.640 242.270 ;
        RECT 2937.860 239.490 2939.040 240.670 ;
        RECT 2939.460 239.490 2940.640 240.670 ;
        RECT 2937.860 61.090 2939.040 62.270 ;
        RECT 2939.460 61.090 2940.640 62.270 ;
        RECT 2937.860 59.490 2939.040 60.670 ;
        RECT 2939.460 59.490 2940.640 60.670 ;
        RECT 2937.860 -14.060 2939.040 -12.880 ;
        RECT 2939.460 -14.060 2940.640 -12.880 ;
        RECT 2937.860 -15.660 2939.040 -14.480 ;
        RECT 2939.460 -15.660 2940.640 -14.480 ;
      LAYER met5 ;
        RECT -21.180 3532.400 2940.800 3535.500 ;
        RECT -45.180 3479.330 2964.800 3482.430 ;
        RECT -45.180 3299.330 2964.800 3302.430 ;
        RECT -45.180 3119.330 2964.800 3122.430 ;
        RECT -45.180 2939.330 2964.800 2942.430 ;
        RECT -45.180 2759.330 2964.800 2762.430 ;
        RECT -45.180 2579.330 2964.800 2582.430 ;
        RECT -45.180 2399.330 2964.800 2402.430 ;
        RECT -45.180 2219.330 2964.800 2222.430 ;
        RECT -45.180 2039.330 2964.800 2042.430 ;
        RECT -45.180 1859.330 2964.800 1862.430 ;
        RECT -45.180 1679.330 2964.800 1682.430 ;
        RECT -45.180 1499.330 2964.800 1502.430 ;
        RECT -45.180 1319.330 2964.800 1322.430 ;
        RECT -45.180 1139.330 2964.800 1142.430 ;
        RECT -45.180 959.330 2964.800 962.430 ;
        RECT -45.180 779.330 2964.800 782.430 ;
        RECT -45.180 599.330 2964.800 602.430 ;
        RECT -45.180 419.330 2964.800 422.430 ;
        RECT -45.180 239.330 2964.800 242.430 ;
        RECT -45.180 59.330 2964.800 62.430 ;
        RECT -21.180 -15.820 2940.800 -12.720 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -30.780 -25.420 -27.680 3545.100 ;
        RECT 98.970 -39.820 102.070 3559.500 ;
        RECT 278.970 -39.820 282.070 3559.500 ;
        RECT 458.970 760.000 462.070 3559.500 ;
        RECT 638.970 760.000 642.070 3559.500 ;
        RECT 458.970 -39.820 462.070 490.000 ;
        RECT 638.970 -39.820 642.070 490.000 ;
        RECT 818.970 -39.820 822.070 3559.500 ;
        RECT 998.970 -39.820 1002.070 3559.500 ;
        RECT 1178.970 -39.820 1182.070 3559.500 ;
        RECT 1358.970 -39.820 1362.070 3559.500 ;
        RECT 1538.970 -39.820 1542.070 3559.500 ;
        RECT 1718.970 -39.820 1722.070 3559.500 ;
        RECT 1898.970 -39.820 1902.070 3559.500 ;
        RECT 2078.970 -39.820 2082.070 3559.500 ;
        RECT 2258.970 -39.820 2262.070 3559.500 ;
        RECT 2438.970 -39.820 2442.070 3559.500 ;
        RECT 2618.970 -39.820 2622.070 3559.500 ;
        RECT 2798.970 -39.820 2802.070 3559.500 ;
        RECT 2947.300 -25.420 2950.400 3545.100 ;
      LAYER via4 ;
        RECT -30.620 3543.760 -29.440 3544.940 ;
        RECT -29.020 3543.760 -27.840 3544.940 ;
        RECT -30.620 3542.160 -29.440 3543.340 ;
        RECT -29.020 3542.160 -27.840 3543.340 ;
        RECT -30.620 3346.090 -29.440 3347.270 ;
        RECT -29.020 3346.090 -27.840 3347.270 ;
        RECT -30.620 3344.490 -29.440 3345.670 ;
        RECT -29.020 3344.490 -27.840 3345.670 ;
        RECT -30.620 3166.090 -29.440 3167.270 ;
        RECT -29.020 3166.090 -27.840 3167.270 ;
        RECT -30.620 3164.490 -29.440 3165.670 ;
        RECT -29.020 3164.490 -27.840 3165.670 ;
        RECT -30.620 2986.090 -29.440 2987.270 ;
        RECT -29.020 2986.090 -27.840 2987.270 ;
        RECT -30.620 2984.490 -29.440 2985.670 ;
        RECT -29.020 2984.490 -27.840 2985.670 ;
        RECT -30.620 2806.090 -29.440 2807.270 ;
        RECT -29.020 2806.090 -27.840 2807.270 ;
        RECT -30.620 2804.490 -29.440 2805.670 ;
        RECT -29.020 2804.490 -27.840 2805.670 ;
        RECT -30.620 2626.090 -29.440 2627.270 ;
        RECT -29.020 2626.090 -27.840 2627.270 ;
        RECT -30.620 2624.490 -29.440 2625.670 ;
        RECT -29.020 2624.490 -27.840 2625.670 ;
        RECT -30.620 2446.090 -29.440 2447.270 ;
        RECT -29.020 2446.090 -27.840 2447.270 ;
        RECT -30.620 2444.490 -29.440 2445.670 ;
        RECT -29.020 2444.490 -27.840 2445.670 ;
        RECT -30.620 2266.090 -29.440 2267.270 ;
        RECT -29.020 2266.090 -27.840 2267.270 ;
        RECT -30.620 2264.490 -29.440 2265.670 ;
        RECT -29.020 2264.490 -27.840 2265.670 ;
        RECT -30.620 2086.090 -29.440 2087.270 ;
        RECT -29.020 2086.090 -27.840 2087.270 ;
        RECT -30.620 2084.490 -29.440 2085.670 ;
        RECT -29.020 2084.490 -27.840 2085.670 ;
        RECT -30.620 1906.090 -29.440 1907.270 ;
        RECT -29.020 1906.090 -27.840 1907.270 ;
        RECT -30.620 1904.490 -29.440 1905.670 ;
        RECT -29.020 1904.490 -27.840 1905.670 ;
        RECT -30.620 1726.090 -29.440 1727.270 ;
        RECT -29.020 1726.090 -27.840 1727.270 ;
        RECT -30.620 1724.490 -29.440 1725.670 ;
        RECT -29.020 1724.490 -27.840 1725.670 ;
        RECT -30.620 1546.090 -29.440 1547.270 ;
        RECT -29.020 1546.090 -27.840 1547.270 ;
        RECT -30.620 1544.490 -29.440 1545.670 ;
        RECT -29.020 1544.490 -27.840 1545.670 ;
        RECT -30.620 1366.090 -29.440 1367.270 ;
        RECT -29.020 1366.090 -27.840 1367.270 ;
        RECT -30.620 1364.490 -29.440 1365.670 ;
        RECT -29.020 1364.490 -27.840 1365.670 ;
        RECT -30.620 1186.090 -29.440 1187.270 ;
        RECT -29.020 1186.090 -27.840 1187.270 ;
        RECT -30.620 1184.490 -29.440 1185.670 ;
        RECT -29.020 1184.490 -27.840 1185.670 ;
        RECT -30.620 1006.090 -29.440 1007.270 ;
        RECT -29.020 1006.090 -27.840 1007.270 ;
        RECT -30.620 1004.490 -29.440 1005.670 ;
        RECT -29.020 1004.490 -27.840 1005.670 ;
        RECT -30.620 826.090 -29.440 827.270 ;
        RECT -29.020 826.090 -27.840 827.270 ;
        RECT -30.620 824.490 -29.440 825.670 ;
        RECT -29.020 824.490 -27.840 825.670 ;
        RECT -30.620 646.090 -29.440 647.270 ;
        RECT -29.020 646.090 -27.840 647.270 ;
        RECT -30.620 644.490 -29.440 645.670 ;
        RECT -29.020 644.490 -27.840 645.670 ;
        RECT -30.620 466.090 -29.440 467.270 ;
        RECT -29.020 466.090 -27.840 467.270 ;
        RECT -30.620 464.490 -29.440 465.670 ;
        RECT -29.020 464.490 -27.840 465.670 ;
        RECT -30.620 286.090 -29.440 287.270 ;
        RECT -29.020 286.090 -27.840 287.270 ;
        RECT -30.620 284.490 -29.440 285.670 ;
        RECT -29.020 284.490 -27.840 285.670 ;
        RECT -30.620 106.090 -29.440 107.270 ;
        RECT -29.020 106.090 -27.840 107.270 ;
        RECT -30.620 104.490 -29.440 105.670 ;
        RECT -29.020 104.490 -27.840 105.670 ;
        RECT -30.620 -23.660 -29.440 -22.480 ;
        RECT -29.020 -23.660 -27.840 -22.480 ;
        RECT -30.620 -25.260 -29.440 -24.080 ;
        RECT -29.020 -25.260 -27.840 -24.080 ;
        RECT 99.130 3543.760 100.310 3544.940 ;
        RECT 100.730 3543.760 101.910 3544.940 ;
        RECT 99.130 3542.160 100.310 3543.340 ;
        RECT 100.730 3542.160 101.910 3543.340 ;
        RECT 99.130 3346.090 100.310 3347.270 ;
        RECT 100.730 3346.090 101.910 3347.270 ;
        RECT 99.130 3344.490 100.310 3345.670 ;
        RECT 100.730 3344.490 101.910 3345.670 ;
        RECT 99.130 3166.090 100.310 3167.270 ;
        RECT 100.730 3166.090 101.910 3167.270 ;
        RECT 99.130 3164.490 100.310 3165.670 ;
        RECT 100.730 3164.490 101.910 3165.670 ;
        RECT 99.130 2986.090 100.310 2987.270 ;
        RECT 100.730 2986.090 101.910 2987.270 ;
        RECT 99.130 2984.490 100.310 2985.670 ;
        RECT 100.730 2984.490 101.910 2985.670 ;
        RECT 99.130 2806.090 100.310 2807.270 ;
        RECT 100.730 2806.090 101.910 2807.270 ;
        RECT 99.130 2804.490 100.310 2805.670 ;
        RECT 100.730 2804.490 101.910 2805.670 ;
        RECT 99.130 2626.090 100.310 2627.270 ;
        RECT 100.730 2626.090 101.910 2627.270 ;
        RECT 99.130 2624.490 100.310 2625.670 ;
        RECT 100.730 2624.490 101.910 2625.670 ;
        RECT 99.130 2446.090 100.310 2447.270 ;
        RECT 100.730 2446.090 101.910 2447.270 ;
        RECT 99.130 2444.490 100.310 2445.670 ;
        RECT 100.730 2444.490 101.910 2445.670 ;
        RECT 99.130 2266.090 100.310 2267.270 ;
        RECT 100.730 2266.090 101.910 2267.270 ;
        RECT 99.130 2264.490 100.310 2265.670 ;
        RECT 100.730 2264.490 101.910 2265.670 ;
        RECT 99.130 2086.090 100.310 2087.270 ;
        RECT 100.730 2086.090 101.910 2087.270 ;
        RECT 99.130 2084.490 100.310 2085.670 ;
        RECT 100.730 2084.490 101.910 2085.670 ;
        RECT 99.130 1906.090 100.310 1907.270 ;
        RECT 100.730 1906.090 101.910 1907.270 ;
        RECT 99.130 1904.490 100.310 1905.670 ;
        RECT 100.730 1904.490 101.910 1905.670 ;
        RECT 99.130 1726.090 100.310 1727.270 ;
        RECT 100.730 1726.090 101.910 1727.270 ;
        RECT 99.130 1724.490 100.310 1725.670 ;
        RECT 100.730 1724.490 101.910 1725.670 ;
        RECT 99.130 1546.090 100.310 1547.270 ;
        RECT 100.730 1546.090 101.910 1547.270 ;
        RECT 99.130 1544.490 100.310 1545.670 ;
        RECT 100.730 1544.490 101.910 1545.670 ;
        RECT 99.130 1366.090 100.310 1367.270 ;
        RECT 100.730 1366.090 101.910 1367.270 ;
        RECT 99.130 1364.490 100.310 1365.670 ;
        RECT 100.730 1364.490 101.910 1365.670 ;
        RECT 99.130 1186.090 100.310 1187.270 ;
        RECT 100.730 1186.090 101.910 1187.270 ;
        RECT 99.130 1184.490 100.310 1185.670 ;
        RECT 100.730 1184.490 101.910 1185.670 ;
        RECT 99.130 1006.090 100.310 1007.270 ;
        RECT 100.730 1006.090 101.910 1007.270 ;
        RECT 99.130 1004.490 100.310 1005.670 ;
        RECT 100.730 1004.490 101.910 1005.670 ;
        RECT 99.130 826.090 100.310 827.270 ;
        RECT 100.730 826.090 101.910 827.270 ;
        RECT 99.130 824.490 100.310 825.670 ;
        RECT 100.730 824.490 101.910 825.670 ;
        RECT 99.130 646.090 100.310 647.270 ;
        RECT 100.730 646.090 101.910 647.270 ;
        RECT 99.130 644.490 100.310 645.670 ;
        RECT 100.730 644.490 101.910 645.670 ;
        RECT 99.130 466.090 100.310 467.270 ;
        RECT 100.730 466.090 101.910 467.270 ;
        RECT 99.130 464.490 100.310 465.670 ;
        RECT 100.730 464.490 101.910 465.670 ;
        RECT 99.130 286.090 100.310 287.270 ;
        RECT 100.730 286.090 101.910 287.270 ;
        RECT 99.130 284.490 100.310 285.670 ;
        RECT 100.730 284.490 101.910 285.670 ;
        RECT 99.130 106.090 100.310 107.270 ;
        RECT 100.730 106.090 101.910 107.270 ;
        RECT 99.130 104.490 100.310 105.670 ;
        RECT 100.730 104.490 101.910 105.670 ;
        RECT 99.130 -23.660 100.310 -22.480 ;
        RECT 100.730 -23.660 101.910 -22.480 ;
        RECT 99.130 -25.260 100.310 -24.080 ;
        RECT 100.730 -25.260 101.910 -24.080 ;
        RECT 279.130 3543.760 280.310 3544.940 ;
        RECT 280.730 3543.760 281.910 3544.940 ;
        RECT 279.130 3542.160 280.310 3543.340 ;
        RECT 280.730 3542.160 281.910 3543.340 ;
        RECT 279.130 3346.090 280.310 3347.270 ;
        RECT 280.730 3346.090 281.910 3347.270 ;
        RECT 279.130 3344.490 280.310 3345.670 ;
        RECT 280.730 3344.490 281.910 3345.670 ;
        RECT 279.130 3166.090 280.310 3167.270 ;
        RECT 280.730 3166.090 281.910 3167.270 ;
        RECT 279.130 3164.490 280.310 3165.670 ;
        RECT 280.730 3164.490 281.910 3165.670 ;
        RECT 279.130 2986.090 280.310 2987.270 ;
        RECT 280.730 2986.090 281.910 2987.270 ;
        RECT 279.130 2984.490 280.310 2985.670 ;
        RECT 280.730 2984.490 281.910 2985.670 ;
        RECT 279.130 2806.090 280.310 2807.270 ;
        RECT 280.730 2806.090 281.910 2807.270 ;
        RECT 279.130 2804.490 280.310 2805.670 ;
        RECT 280.730 2804.490 281.910 2805.670 ;
        RECT 279.130 2626.090 280.310 2627.270 ;
        RECT 280.730 2626.090 281.910 2627.270 ;
        RECT 279.130 2624.490 280.310 2625.670 ;
        RECT 280.730 2624.490 281.910 2625.670 ;
        RECT 279.130 2446.090 280.310 2447.270 ;
        RECT 280.730 2446.090 281.910 2447.270 ;
        RECT 279.130 2444.490 280.310 2445.670 ;
        RECT 280.730 2444.490 281.910 2445.670 ;
        RECT 279.130 2266.090 280.310 2267.270 ;
        RECT 280.730 2266.090 281.910 2267.270 ;
        RECT 279.130 2264.490 280.310 2265.670 ;
        RECT 280.730 2264.490 281.910 2265.670 ;
        RECT 279.130 2086.090 280.310 2087.270 ;
        RECT 280.730 2086.090 281.910 2087.270 ;
        RECT 279.130 2084.490 280.310 2085.670 ;
        RECT 280.730 2084.490 281.910 2085.670 ;
        RECT 279.130 1906.090 280.310 1907.270 ;
        RECT 280.730 1906.090 281.910 1907.270 ;
        RECT 279.130 1904.490 280.310 1905.670 ;
        RECT 280.730 1904.490 281.910 1905.670 ;
        RECT 279.130 1726.090 280.310 1727.270 ;
        RECT 280.730 1726.090 281.910 1727.270 ;
        RECT 279.130 1724.490 280.310 1725.670 ;
        RECT 280.730 1724.490 281.910 1725.670 ;
        RECT 279.130 1546.090 280.310 1547.270 ;
        RECT 280.730 1546.090 281.910 1547.270 ;
        RECT 279.130 1544.490 280.310 1545.670 ;
        RECT 280.730 1544.490 281.910 1545.670 ;
        RECT 279.130 1366.090 280.310 1367.270 ;
        RECT 280.730 1366.090 281.910 1367.270 ;
        RECT 279.130 1364.490 280.310 1365.670 ;
        RECT 280.730 1364.490 281.910 1365.670 ;
        RECT 279.130 1186.090 280.310 1187.270 ;
        RECT 280.730 1186.090 281.910 1187.270 ;
        RECT 279.130 1184.490 280.310 1185.670 ;
        RECT 280.730 1184.490 281.910 1185.670 ;
        RECT 279.130 1006.090 280.310 1007.270 ;
        RECT 280.730 1006.090 281.910 1007.270 ;
        RECT 279.130 1004.490 280.310 1005.670 ;
        RECT 280.730 1004.490 281.910 1005.670 ;
        RECT 279.130 826.090 280.310 827.270 ;
        RECT 280.730 826.090 281.910 827.270 ;
        RECT 279.130 824.490 280.310 825.670 ;
        RECT 280.730 824.490 281.910 825.670 ;
        RECT 459.130 3543.760 460.310 3544.940 ;
        RECT 460.730 3543.760 461.910 3544.940 ;
        RECT 459.130 3542.160 460.310 3543.340 ;
        RECT 460.730 3542.160 461.910 3543.340 ;
        RECT 459.130 3346.090 460.310 3347.270 ;
        RECT 460.730 3346.090 461.910 3347.270 ;
        RECT 459.130 3344.490 460.310 3345.670 ;
        RECT 460.730 3344.490 461.910 3345.670 ;
        RECT 459.130 3166.090 460.310 3167.270 ;
        RECT 460.730 3166.090 461.910 3167.270 ;
        RECT 459.130 3164.490 460.310 3165.670 ;
        RECT 460.730 3164.490 461.910 3165.670 ;
        RECT 459.130 2986.090 460.310 2987.270 ;
        RECT 460.730 2986.090 461.910 2987.270 ;
        RECT 459.130 2984.490 460.310 2985.670 ;
        RECT 460.730 2984.490 461.910 2985.670 ;
        RECT 459.130 2806.090 460.310 2807.270 ;
        RECT 460.730 2806.090 461.910 2807.270 ;
        RECT 459.130 2804.490 460.310 2805.670 ;
        RECT 460.730 2804.490 461.910 2805.670 ;
        RECT 459.130 2626.090 460.310 2627.270 ;
        RECT 460.730 2626.090 461.910 2627.270 ;
        RECT 459.130 2624.490 460.310 2625.670 ;
        RECT 460.730 2624.490 461.910 2625.670 ;
        RECT 459.130 2446.090 460.310 2447.270 ;
        RECT 460.730 2446.090 461.910 2447.270 ;
        RECT 459.130 2444.490 460.310 2445.670 ;
        RECT 460.730 2444.490 461.910 2445.670 ;
        RECT 459.130 2266.090 460.310 2267.270 ;
        RECT 460.730 2266.090 461.910 2267.270 ;
        RECT 459.130 2264.490 460.310 2265.670 ;
        RECT 460.730 2264.490 461.910 2265.670 ;
        RECT 459.130 2086.090 460.310 2087.270 ;
        RECT 460.730 2086.090 461.910 2087.270 ;
        RECT 459.130 2084.490 460.310 2085.670 ;
        RECT 460.730 2084.490 461.910 2085.670 ;
        RECT 459.130 1906.090 460.310 1907.270 ;
        RECT 460.730 1906.090 461.910 1907.270 ;
        RECT 459.130 1904.490 460.310 1905.670 ;
        RECT 460.730 1904.490 461.910 1905.670 ;
        RECT 459.130 1726.090 460.310 1727.270 ;
        RECT 460.730 1726.090 461.910 1727.270 ;
        RECT 459.130 1724.490 460.310 1725.670 ;
        RECT 460.730 1724.490 461.910 1725.670 ;
        RECT 459.130 1546.090 460.310 1547.270 ;
        RECT 460.730 1546.090 461.910 1547.270 ;
        RECT 459.130 1544.490 460.310 1545.670 ;
        RECT 460.730 1544.490 461.910 1545.670 ;
        RECT 459.130 1366.090 460.310 1367.270 ;
        RECT 460.730 1366.090 461.910 1367.270 ;
        RECT 459.130 1364.490 460.310 1365.670 ;
        RECT 460.730 1364.490 461.910 1365.670 ;
        RECT 459.130 1186.090 460.310 1187.270 ;
        RECT 460.730 1186.090 461.910 1187.270 ;
        RECT 459.130 1184.490 460.310 1185.670 ;
        RECT 460.730 1184.490 461.910 1185.670 ;
        RECT 459.130 1006.090 460.310 1007.270 ;
        RECT 460.730 1006.090 461.910 1007.270 ;
        RECT 459.130 1004.490 460.310 1005.670 ;
        RECT 460.730 1004.490 461.910 1005.670 ;
        RECT 459.130 826.090 460.310 827.270 ;
        RECT 460.730 826.090 461.910 827.270 ;
        RECT 459.130 824.490 460.310 825.670 ;
        RECT 460.730 824.490 461.910 825.670 ;
        RECT 639.130 3543.760 640.310 3544.940 ;
        RECT 640.730 3543.760 641.910 3544.940 ;
        RECT 639.130 3542.160 640.310 3543.340 ;
        RECT 640.730 3542.160 641.910 3543.340 ;
        RECT 639.130 3346.090 640.310 3347.270 ;
        RECT 640.730 3346.090 641.910 3347.270 ;
        RECT 639.130 3344.490 640.310 3345.670 ;
        RECT 640.730 3344.490 641.910 3345.670 ;
        RECT 639.130 3166.090 640.310 3167.270 ;
        RECT 640.730 3166.090 641.910 3167.270 ;
        RECT 639.130 3164.490 640.310 3165.670 ;
        RECT 640.730 3164.490 641.910 3165.670 ;
        RECT 639.130 2986.090 640.310 2987.270 ;
        RECT 640.730 2986.090 641.910 2987.270 ;
        RECT 639.130 2984.490 640.310 2985.670 ;
        RECT 640.730 2984.490 641.910 2985.670 ;
        RECT 639.130 2806.090 640.310 2807.270 ;
        RECT 640.730 2806.090 641.910 2807.270 ;
        RECT 639.130 2804.490 640.310 2805.670 ;
        RECT 640.730 2804.490 641.910 2805.670 ;
        RECT 639.130 2626.090 640.310 2627.270 ;
        RECT 640.730 2626.090 641.910 2627.270 ;
        RECT 639.130 2624.490 640.310 2625.670 ;
        RECT 640.730 2624.490 641.910 2625.670 ;
        RECT 639.130 2446.090 640.310 2447.270 ;
        RECT 640.730 2446.090 641.910 2447.270 ;
        RECT 639.130 2444.490 640.310 2445.670 ;
        RECT 640.730 2444.490 641.910 2445.670 ;
        RECT 639.130 2266.090 640.310 2267.270 ;
        RECT 640.730 2266.090 641.910 2267.270 ;
        RECT 639.130 2264.490 640.310 2265.670 ;
        RECT 640.730 2264.490 641.910 2265.670 ;
        RECT 639.130 2086.090 640.310 2087.270 ;
        RECT 640.730 2086.090 641.910 2087.270 ;
        RECT 639.130 2084.490 640.310 2085.670 ;
        RECT 640.730 2084.490 641.910 2085.670 ;
        RECT 639.130 1906.090 640.310 1907.270 ;
        RECT 640.730 1906.090 641.910 1907.270 ;
        RECT 639.130 1904.490 640.310 1905.670 ;
        RECT 640.730 1904.490 641.910 1905.670 ;
        RECT 639.130 1726.090 640.310 1727.270 ;
        RECT 640.730 1726.090 641.910 1727.270 ;
        RECT 639.130 1724.490 640.310 1725.670 ;
        RECT 640.730 1724.490 641.910 1725.670 ;
        RECT 639.130 1546.090 640.310 1547.270 ;
        RECT 640.730 1546.090 641.910 1547.270 ;
        RECT 639.130 1544.490 640.310 1545.670 ;
        RECT 640.730 1544.490 641.910 1545.670 ;
        RECT 639.130 1366.090 640.310 1367.270 ;
        RECT 640.730 1366.090 641.910 1367.270 ;
        RECT 639.130 1364.490 640.310 1365.670 ;
        RECT 640.730 1364.490 641.910 1365.670 ;
        RECT 639.130 1186.090 640.310 1187.270 ;
        RECT 640.730 1186.090 641.910 1187.270 ;
        RECT 639.130 1184.490 640.310 1185.670 ;
        RECT 640.730 1184.490 641.910 1185.670 ;
        RECT 639.130 1006.090 640.310 1007.270 ;
        RECT 640.730 1006.090 641.910 1007.270 ;
        RECT 639.130 1004.490 640.310 1005.670 ;
        RECT 640.730 1004.490 641.910 1005.670 ;
        RECT 639.130 826.090 640.310 827.270 ;
        RECT 640.730 826.090 641.910 827.270 ;
        RECT 639.130 824.490 640.310 825.670 ;
        RECT 640.730 824.490 641.910 825.670 ;
        RECT 819.130 3543.760 820.310 3544.940 ;
        RECT 820.730 3543.760 821.910 3544.940 ;
        RECT 819.130 3542.160 820.310 3543.340 ;
        RECT 820.730 3542.160 821.910 3543.340 ;
        RECT 819.130 3346.090 820.310 3347.270 ;
        RECT 820.730 3346.090 821.910 3347.270 ;
        RECT 819.130 3344.490 820.310 3345.670 ;
        RECT 820.730 3344.490 821.910 3345.670 ;
        RECT 819.130 3166.090 820.310 3167.270 ;
        RECT 820.730 3166.090 821.910 3167.270 ;
        RECT 819.130 3164.490 820.310 3165.670 ;
        RECT 820.730 3164.490 821.910 3165.670 ;
        RECT 819.130 2986.090 820.310 2987.270 ;
        RECT 820.730 2986.090 821.910 2987.270 ;
        RECT 819.130 2984.490 820.310 2985.670 ;
        RECT 820.730 2984.490 821.910 2985.670 ;
        RECT 819.130 2806.090 820.310 2807.270 ;
        RECT 820.730 2806.090 821.910 2807.270 ;
        RECT 819.130 2804.490 820.310 2805.670 ;
        RECT 820.730 2804.490 821.910 2805.670 ;
        RECT 819.130 2626.090 820.310 2627.270 ;
        RECT 820.730 2626.090 821.910 2627.270 ;
        RECT 819.130 2624.490 820.310 2625.670 ;
        RECT 820.730 2624.490 821.910 2625.670 ;
        RECT 819.130 2446.090 820.310 2447.270 ;
        RECT 820.730 2446.090 821.910 2447.270 ;
        RECT 819.130 2444.490 820.310 2445.670 ;
        RECT 820.730 2444.490 821.910 2445.670 ;
        RECT 819.130 2266.090 820.310 2267.270 ;
        RECT 820.730 2266.090 821.910 2267.270 ;
        RECT 819.130 2264.490 820.310 2265.670 ;
        RECT 820.730 2264.490 821.910 2265.670 ;
        RECT 819.130 2086.090 820.310 2087.270 ;
        RECT 820.730 2086.090 821.910 2087.270 ;
        RECT 819.130 2084.490 820.310 2085.670 ;
        RECT 820.730 2084.490 821.910 2085.670 ;
        RECT 819.130 1906.090 820.310 1907.270 ;
        RECT 820.730 1906.090 821.910 1907.270 ;
        RECT 819.130 1904.490 820.310 1905.670 ;
        RECT 820.730 1904.490 821.910 1905.670 ;
        RECT 819.130 1726.090 820.310 1727.270 ;
        RECT 820.730 1726.090 821.910 1727.270 ;
        RECT 819.130 1724.490 820.310 1725.670 ;
        RECT 820.730 1724.490 821.910 1725.670 ;
        RECT 819.130 1546.090 820.310 1547.270 ;
        RECT 820.730 1546.090 821.910 1547.270 ;
        RECT 819.130 1544.490 820.310 1545.670 ;
        RECT 820.730 1544.490 821.910 1545.670 ;
        RECT 819.130 1366.090 820.310 1367.270 ;
        RECT 820.730 1366.090 821.910 1367.270 ;
        RECT 819.130 1364.490 820.310 1365.670 ;
        RECT 820.730 1364.490 821.910 1365.670 ;
        RECT 819.130 1186.090 820.310 1187.270 ;
        RECT 820.730 1186.090 821.910 1187.270 ;
        RECT 819.130 1184.490 820.310 1185.670 ;
        RECT 820.730 1184.490 821.910 1185.670 ;
        RECT 819.130 1006.090 820.310 1007.270 ;
        RECT 820.730 1006.090 821.910 1007.270 ;
        RECT 819.130 1004.490 820.310 1005.670 ;
        RECT 820.730 1004.490 821.910 1005.670 ;
        RECT 819.130 826.090 820.310 827.270 ;
        RECT 820.730 826.090 821.910 827.270 ;
        RECT 819.130 824.490 820.310 825.670 ;
        RECT 820.730 824.490 821.910 825.670 ;
        RECT 279.130 646.090 280.310 647.270 ;
        RECT 280.730 646.090 281.910 647.270 ;
        RECT 279.130 644.490 280.310 645.670 ;
        RECT 280.730 644.490 281.910 645.670 ;
        RECT 819.130 646.090 820.310 647.270 ;
        RECT 820.730 646.090 821.910 647.270 ;
        RECT 819.130 644.490 820.310 645.670 ;
        RECT 820.730 644.490 821.910 645.670 ;
        RECT 279.130 466.090 280.310 467.270 ;
        RECT 280.730 466.090 281.910 467.270 ;
        RECT 279.130 464.490 280.310 465.670 ;
        RECT 280.730 464.490 281.910 465.670 ;
        RECT 279.130 286.090 280.310 287.270 ;
        RECT 280.730 286.090 281.910 287.270 ;
        RECT 279.130 284.490 280.310 285.670 ;
        RECT 280.730 284.490 281.910 285.670 ;
        RECT 279.130 106.090 280.310 107.270 ;
        RECT 280.730 106.090 281.910 107.270 ;
        RECT 279.130 104.490 280.310 105.670 ;
        RECT 280.730 104.490 281.910 105.670 ;
        RECT 279.130 -23.660 280.310 -22.480 ;
        RECT 280.730 -23.660 281.910 -22.480 ;
        RECT 279.130 -25.260 280.310 -24.080 ;
        RECT 280.730 -25.260 281.910 -24.080 ;
        RECT 459.130 466.090 460.310 467.270 ;
        RECT 460.730 466.090 461.910 467.270 ;
        RECT 459.130 464.490 460.310 465.670 ;
        RECT 460.730 464.490 461.910 465.670 ;
        RECT 459.130 286.090 460.310 287.270 ;
        RECT 460.730 286.090 461.910 287.270 ;
        RECT 459.130 284.490 460.310 285.670 ;
        RECT 460.730 284.490 461.910 285.670 ;
        RECT 459.130 106.090 460.310 107.270 ;
        RECT 460.730 106.090 461.910 107.270 ;
        RECT 459.130 104.490 460.310 105.670 ;
        RECT 460.730 104.490 461.910 105.670 ;
        RECT 459.130 -23.660 460.310 -22.480 ;
        RECT 460.730 -23.660 461.910 -22.480 ;
        RECT 459.130 -25.260 460.310 -24.080 ;
        RECT 460.730 -25.260 461.910 -24.080 ;
        RECT 639.130 466.090 640.310 467.270 ;
        RECT 640.730 466.090 641.910 467.270 ;
        RECT 639.130 464.490 640.310 465.670 ;
        RECT 640.730 464.490 641.910 465.670 ;
        RECT 639.130 286.090 640.310 287.270 ;
        RECT 640.730 286.090 641.910 287.270 ;
        RECT 639.130 284.490 640.310 285.670 ;
        RECT 640.730 284.490 641.910 285.670 ;
        RECT 639.130 106.090 640.310 107.270 ;
        RECT 640.730 106.090 641.910 107.270 ;
        RECT 639.130 104.490 640.310 105.670 ;
        RECT 640.730 104.490 641.910 105.670 ;
        RECT 639.130 -23.660 640.310 -22.480 ;
        RECT 640.730 -23.660 641.910 -22.480 ;
        RECT 639.130 -25.260 640.310 -24.080 ;
        RECT 640.730 -25.260 641.910 -24.080 ;
        RECT 819.130 466.090 820.310 467.270 ;
        RECT 820.730 466.090 821.910 467.270 ;
        RECT 819.130 464.490 820.310 465.670 ;
        RECT 820.730 464.490 821.910 465.670 ;
        RECT 819.130 286.090 820.310 287.270 ;
        RECT 820.730 286.090 821.910 287.270 ;
        RECT 819.130 284.490 820.310 285.670 ;
        RECT 820.730 284.490 821.910 285.670 ;
        RECT 819.130 106.090 820.310 107.270 ;
        RECT 820.730 106.090 821.910 107.270 ;
        RECT 819.130 104.490 820.310 105.670 ;
        RECT 820.730 104.490 821.910 105.670 ;
        RECT 819.130 -23.660 820.310 -22.480 ;
        RECT 820.730 -23.660 821.910 -22.480 ;
        RECT 819.130 -25.260 820.310 -24.080 ;
        RECT 820.730 -25.260 821.910 -24.080 ;
        RECT 999.130 3543.760 1000.310 3544.940 ;
        RECT 1000.730 3543.760 1001.910 3544.940 ;
        RECT 999.130 3542.160 1000.310 3543.340 ;
        RECT 1000.730 3542.160 1001.910 3543.340 ;
        RECT 999.130 3346.090 1000.310 3347.270 ;
        RECT 1000.730 3346.090 1001.910 3347.270 ;
        RECT 999.130 3344.490 1000.310 3345.670 ;
        RECT 1000.730 3344.490 1001.910 3345.670 ;
        RECT 999.130 3166.090 1000.310 3167.270 ;
        RECT 1000.730 3166.090 1001.910 3167.270 ;
        RECT 999.130 3164.490 1000.310 3165.670 ;
        RECT 1000.730 3164.490 1001.910 3165.670 ;
        RECT 999.130 2986.090 1000.310 2987.270 ;
        RECT 1000.730 2986.090 1001.910 2987.270 ;
        RECT 999.130 2984.490 1000.310 2985.670 ;
        RECT 1000.730 2984.490 1001.910 2985.670 ;
        RECT 999.130 2806.090 1000.310 2807.270 ;
        RECT 1000.730 2806.090 1001.910 2807.270 ;
        RECT 999.130 2804.490 1000.310 2805.670 ;
        RECT 1000.730 2804.490 1001.910 2805.670 ;
        RECT 999.130 2626.090 1000.310 2627.270 ;
        RECT 1000.730 2626.090 1001.910 2627.270 ;
        RECT 999.130 2624.490 1000.310 2625.670 ;
        RECT 1000.730 2624.490 1001.910 2625.670 ;
        RECT 999.130 2446.090 1000.310 2447.270 ;
        RECT 1000.730 2446.090 1001.910 2447.270 ;
        RECT 999.130 2444.490 1000.310 2445.670 ;
        RECT 1000.730 2444.490 1001.910 2445.670 ;
        RECT 999.130 2266.090 1000.310 2267.270 ;
        RECT 1000.730 2266.090 1001.910 2267.270 ;
        RECT 999.130 2264.490 1000.310 2265.670 ;
        RECT 1000.730 2264.490 1001.910 2265.670 ;
        RECT 999.130 2086.090 1000.310 2087.270 ;
        RECT 1000.730 2086.090 1001.910 2087.270 ;
        RECT 999.130 2084.490 1000.310 2085.670 ;
        RECT 1000.730 2084.490 1001.910 2085.670 ;
        RECT 999.130 1906.090 1000.310 1907.270 ;
        RECT 1000.730 1906.090 1001.910 1907.270 ;
        RECT 999.130 1904.490 1000.310 1905.670 ;
        RECT 1000.730 1904.490 1001.910 1905.670 ;
        RECT 999.130 1726.090 1000.310 1727.270 ;
        RECT 1000.730 1726.090 1001.910 1727.270 ;
        RECT 999.130 1724.490 1000.310 1725.670 ;
        RECT 1000.730 1724.490 1001.910 1725.670 ;
        RECT 999.130 1546.090 1000.310 1547.270 ;
        RECT 1000.730 1546.090 1001.910 1547.270 ;
        RECT 999.130 1544.490 1000.310 1545.670 ;
        RECT 1000.730 1544.490 1001.910 1545.670 ;
        RECT 999.130 1366.090 1000.310 1367.270 ;
        RECT 1000.730 1366.090 1001.910 1367.270 ;
        RECT 999.130 1364.490 1000.310 1365.670 ;
        RECT 1000.730 1364.490 1001.910 1365.670 ;
        RECT 999.130 1186.090 1000.310 1187.270 ;
        RECT 1000.730 1186.090 1001.910 1187.270 ;
        RECT 999.130 1184.490 1000.310 1185.670 ;
        RECT 1000.730 1184.490 1001.910 1185.670 ;
        RECT 999.130 1006.090 1000.310 1007.270 ;
        RECT 1000.730 1006.090 1001.910 1007.270 ;
        RECT 999.130 1004.490 1000.310 1005.670 ;
        RECT 1000.730 1004.490 1001.910 1005.670 ;
        RECT 999.130 826.090 1000.310 827.270 ;
        RECT 1000.730 826.090 1001.910 827.270 ;
        RECT 999.130 824.490 1000.310 825.670 ;
        RECT 1000.730 824.490 1001.910 825.670 ;
        RECT 999.130 646.090 1000.310 647.270 ;
        RECT 1000.730 646.090 1001.910 647.270 ;
        RECT 999.130 644.490 1000.310 645.670 ;
        RECT 1000.730 644.490 1001.910 645.670 ;
        RECT 999.130 466.090 1000.310 467.270 ;
        RECT 1000.730 466.090 1001.910 467.270 ;
        RECT 999.130 464.490 1000.310 465.670 ;
        RECT 1000.730 464.490 1001.910 465.670 ;
        RECT 999.130 286.090 1000.310 287.270 ;
        RECT 1000.730 286.090 1001.910 287.270 ;
        RECT 999.130 284.490 1000.310 285.670 ;
        RECT 1000.730 284.490 1001.910 285.670 ;
        RECT 999.130 106.090 1000.310 107.270 ;
        RECT 1000.730 106.090 1001.910 107.270 ;
        RECT 999.130 104.490 1000.310 105.670 ;
        RECT 1000.730 104.490 1001.910 105.670 ;
        RECT 999.130 -23.660 1000.310 -22.480 ;
        RECT 1000.730 -23.660 1001.910 -22.480 ;
        RECT 999.130 -25.260 1000.310 -24.080 ;
        RECT 1000.730 -25.260 1001.910 -24.080 ;
        RECT 1179.130 3543.760 1180.310 3544.940 ;
        RECT 1180.730 3543.760 1181.910 3544.940 ;
        RECT 1179.130 3542.160 1180.310 3543.340 ;
        RECT 1180.730 3542.160 1181.910 3543.340 ;
        RECT 1179.130 3346.090 1180.310 3347.270 ;
        RECT 1180.730 3346.090 1181.910 3347.270 ;
        RECT 1179.130 3344.490 1180.310 3345.670 ;
        RECT 1180.730 3344.490 1181.910 3345.670 ;
        RECT 1179.130 3166.090 1180.310 3167.270 ;
        RECT 1180.730 3166.090 1181.910 3167.270 ;
        RECT 1179.130 3164.490 1180.310 3165.670 ;
        RECT 1180.730 3164.490 1181.910 3165.670 ;
        RECT 1179.130 2986.090 1180.310 2987.270 ;
        RECT 1180.730 2986.090 1181.910 2987.270 ;
        RECT 1179.130 2984.490 1180.310 2985.670 ;
        RECT 1180.730 2984.490 1181.910 2985.670 ;
        RECT 1179.130 2806.090 1180.310 2807.270 ;
        RECT 1180.730 2806.090 1181.910 2807.270 ;
        RECT 1179.130 2804.490 1180.310 2805.670 ;
        RECT 1180.730 2804.490 1181.910 2805.670 ;
        RECT 1179.130 2626.090 1180.310 2627.270 ;
        RECT 1180.730 2626.090 1181.910 2627.270 ;
        RECT 1179.130 2624.490 1180.310 2625.670 ;
        RECT 1180.730 2624.490 1181.910 2625.670 ;
        RECT 1179.130 2446.090 1180.310 2447.270 ;
        RECT 1180.730 2446.090 1181.910 2447.270 ;
        RECT 1179.130 2444.490 1180.310 2445.670 ;
        RECT 1180.730 2444.490 1181.910 2445.670 ;
        RECT 1179.130 2266.090 1180.310 2267.270 ;
        RECT 1180.730 2266.090 1181.910 2267.270 ;
        RECT 1179.130 2264.490 1180.310 2265.670 ;
        RECT 1180.730 2264.490 1181.910 2265.670 ;
        RECT 1179.130 2086.090 1180.310 2087.270 ;
        RECT 1180.730 2086.090 1181.910 2087.270 ;
        RECT 1179.130 2084.490 1180.310 2085.670 ;
        RECT 1180.730 2084.490 1181.910 2085.670 ;
        RECT 1179.130 1906.090 1180.310 1907.270 ;
        RECT 1180.730 1906.090 1181.910 1907.270 ;
        RECT 1179.130 1904.490 1180.310 1905.670 ;
        RECT 1180.730 1904.490 1181.910 1905.670 ;
        RECT 1179.130 1726.090 1180.310 1727.270 ;
        RECT 1180.730 1726.090 1181.910 1727.270 ;
        RECT 1179.130 1724.490 1180.310 1725.670 ;
        RECT 1180.730 1724.490 1181.910 1725.670 ;
        RECT 1179.130 1546.090 1180.310 1547.270 ;
        RECT 1180.730 1546.090 1181.910 1547.270 ;
        RECT 1179.130 1544.490 1180.310 1545.670 ;
        RECT 1180.730 1544.490 1181.910 1545.670 ;
        RECT 1179.130 1366.090 1180.310 1367.270 ;
        RECT 1180.730 1366.090 1181.910 1367.270 ;
        RECT 1179.130 1364.490 1180.310 1365.670 ;
        RECT 1180.730 1364.490 1181.910 1365.670 ;
        RECT 1179.130 1186.090 1180.310 1187.270 ;
        RECT 1180.730 1186.090 1181.910 1187.270 ;
        RECT 1179.130 1184.490 1180.310 1185.670 ;
        RECT 1180.730 1184.490 1181.910 1185.670 ;
        RECT 1179.130 1006.090 1180.310 1007.270 ;
        RECT 1180.730 1006.090 1181.910 1007.270 ;
        RECT 1179.130 1004.490 1180.310 1005.670 ;
        RECT 1180.730 1004.490 1181.910 1005.670 ;
        RECT 1179.130 826.090 1180.310 827.270 ;
        RECT 1180.730 826.090 1181.910 827.270 ;
        RECT 1179.130 824.490 1180.310 825.670 ;
        RECT 1180.730 824.490 1181.910 825.670 ;
        RECT 1179.130 646.090 1180.310 647.270 ;
        RECT 1180.730 646.090 1181.910 647.270 ;
        RECT 1179.130 644.490 1180.310 645.670 ;
        RECT 1180.730 644.490 1181.910 645.670 ;
        RECT 1179.130 466.090 1180.310 467.270 ;
        RECT 1180.730 466.090 1181.910 467.270 ;
        RECT 1179.130 464.490 1180.310 465.670 ;
        RECT 1180.730 464.490 1181.910 465.670 ;
        RECT 1179.130 286.090 1180.310 287.270 ;
        RECT 1180.730 286.090 1181.910 287.270 ;
        RECT 1179.130 284.490 1180.310 285.670 ;
        RECT 1180.730 284.490 1181.910 285.670 ;
        RECT 1179.130 106.090 1180.310 107.270 ;
        RECT 1180.730 106.090 1181.910 107.270 ;
        RECT 1179.130 104.490 1180.310 105.670 ;
        RECT 1180.730 104.490 1181.910 105.670 ;
        RECT 1179.130 -23.660 1180.310 -22.480 ;
        RECT 1180.730 -23.660 1181.910 -22.480 ;
        RECT 1179.130 -25.260 1180.310 -24.080 ;
        RECT 1180.730 -25.260 1181.910 -24.080 ;
        RECT 1359.130 3543.760 1360.310 3544.940 ;
        RECT 1360.730 3543.760 1361.910 3544.940 ;
        RECT 1359.130 3542.160 1360.310 3543.340 ;
        RECT 1360.730 3542.160 1361.910 3543.340 ;
        RECT 1359.130 3346.090 1360.310 3347.270 ;
        RECT 1360.730 3346.090 1361.910 3347.270 ;
        RECT 1359.130 3344.490 1360.310 3345.670 ;
        RECT 1360.730 3344.490 1361.910 3345.670 ;
        RECT 1359.130 3166.090 1360.310 3167.270 ;
        RECT 1360.730 3166.090 1361.910 3167.270 ;
        RECT 1359.130 3164.490 1360.310 3165.670 ;
        RECT 1360.730 3164.490 1361.910 3165.670 ;
        RECT 1359.130 2986.090 1360.310 2987.270 ;
        RECT 1360.730 2986.090 1361.910 2987.270 ;
        RECT 1359.130 2984.490 1360.310 2985.670 ;
        RECT 1360.730 2984.490 1361.910 2985.670 ;
        RECT 1359.130 2806.090 1360.310 2807.270 ;
        RECT 1360.730 2806.090 1361.910 2807.270 ;
        RECT 1359.130 2804.490 1360.310 2805.670 ;
        RECT 1360.730 2804.490 1361.910 2805.670 ;
        RECT 1359.130 2626.090 1360.310 2627.270 ;
        RECT 1360.730 2626.090 1361.910 2627.270 ;
        RECT 1359.130 2624.490 1360.310 2625.670 ;
        RECT 1360.730 2624.490 1361.910 2625.670 ;
        RECT 1359.130 2446.090 1360.310 2447.270 ;
        RECT 1360.730 2446.090 1361.910 2447.270 ;
        RECT 1359.130 2444.490 1360.310 2445.670 ;
        RECT 1360.730 2444.490 1361.910 2445.670 ;
        RECT 1359.130 2266.090 1360.310 2267.270 ;
        RECT 1360.730 2266.090 1361.910 2267.270 ;
        RECT 1359.130 2264.490 1360.310 2265.670 ;
        RECT 1360.730 2264.490 1361.910 2265.670 ;
        RECT 1359.130 2086.090 1360.310 2087.270 ;
        RECT 1360.730 2086.090 1361.910 2087.270 ;
        RECT 1359.130 2084.490 1360.310 2085.670 ;
        RECT 1360.730 2084.490 1361.910 2085.670 ;
        RECT 1359.130 1906.090 1360.310 1907.270 ;
        RECT 1360.730 1906.090 1361.910 1907.270 ;
        RECT 1359.130 1904.490 1360.310 1905.670 ;
        RECT 1360.730 1904.490 1361.910 1905.670 ;
        RECT 1359.130 1726.090 1360.310 1727.270 ;
        RECT 1360.730 1726.090 1361.910 1727.270 ;
        RECT 1359.130 1724.490 1360.310 1725.670 ;
        RECT 1360.730 1724.490 1361.910 1725.670 ;
        RECT 1359.130 1546.090 1360.310 1547.270 ;
        RECT 1360.730 1546.090 1361.910 1547.270 ;
        RECT 1359.130 1544.490 1360.310 1545.670 ;
        RECT 1360.730 1544.490 1361.910 1545.670 ;
        RECT 1359.130 1366.090 1360.310 1367.270 ;
        RECT 1360.730 1366.090 1361.910 1367.270 ;
        RECT 1359.130 1364.490 1360.310 1365.670 ;
        RECT 1360.730 1364.490 1361.910 1365.670 ;
        RECT 1359.130 1186.090 1360.310 1187.270 ;
        RECT 1360.730 1186.090 1361.910 1187.270 ;
        RECT 1359.130 1184.490 1360.310 1185.670 ;
        RECT 1360.730 1184.490 1361.910 1185.670 ;
        RECT 1359.130 1006.090 1360.310 1007.270 ;
        RECT 1360.730 1006.090 1361.910 1007.270 ;
        RECT 1359.130 1004.490 1360.310 1005.670 ;
        RECT 1360.730 1004.490 1361.910 1005.670 ;
        RECT 1359.130 826.090 1360.310 827.270 ;
        RECT 1360.730 826.090 1361.910 827.270 ;
        RECT 1359.130 824.490 1360.310 825.670 ;
        RECT 1360.730 824.490 1361.910 825.670 ;
        RECT 1359.130 646.090 1360.310 647.270 ;
        RECT 1360.730 646.090 1361.910 647.270 ;
        RECT 1359.130 644.490 1360.310 645.670 ;
        RECT 1360.730 644.490 1361.910 645.670 ;
        RECT 1359.130 466.090 1360.310 467.270 ;
        RECT 1360.730 466.090 1361.910 467.270 ;
        RECT 1359.130 464.490 1360.310 465.670 ;
        RECT 1360.730 464.490 1361.910 465.670 ;
        RECT 1359.130 286.090 1360.310 287.270 ;
        RECT 1360.730 286.090 1361.910 287.270 ;
        RECT 1359.130 284.490 1360.310 285.670 ;
        RECT 1360.730 284.490 1361.910 285.670 ;
        RECT 1359.130 106.090 1360.310 107.270 ;
        RECT 1360.730 106.090 1361.910 107.270 ;
        RECT 1359.130 104.490 1360.310 105.670 ;
        RECT 1360.730 104.490 1361.910 105.670 ;
        RECT 1359.130 -23.660 1360.310 -22.480 ;
        RECT 1360.730 -23.660 1361.910 -22.480 ;
        RECT 1359.130 -25.260 1360.310 -24.080 ;
        RECT 1360.730 -25.260 1361.910 -24.080 ;
        RECT 1539.130 3543.760 1540.310 3544.940 ;
        RECT 1540.730 3543.760 1541.910 3544.940 ;
        RECT 1539.130 3542.160 1540.310 3543.340 ;
        RECT 1540.730 3542.160 1541.910 3543.340 ;
        RECT 1539.130 3346.090 1540.310 3347.270 ;
        RECT 1540.730 3346.090 1541.910 3347.270 ;
        RECT 1539.130 3344.490 1540.310 3345.670 ;
        RECT 1540.730 3344.490 1541.910 3345.670 ;
        RECT 1539.130 3166.090 1540.310 3167.270 ;
        RECT 1540.730 3166.090 1541.910 3167.270 ;
        RECT 1539.130 3164.490 1540.310 3165.670 ;
        RECT 1540.730 3164.490 1541.910 3165.670 ;
        RECT 1539.130 2986.090 1540.310 2987.270 ;
        RECT 1540.730 2986.090 1541.910 2987.270 ;
        RECT 1539.130 2984.490 1540.310 2985.670 ;
        RECT 1540.730 2984.490 1541.910 2985.670 ;
        RECT 1539.130 2806.090 1540.310 2807.270 ;
        RECT 1540.730 2806.090 1541.910 2807.270 ;
        RECT 1539.130 2804.490 1540.310 2805.670 ;
        RECT 1540.730 2804.490 1541.910 2805.670 ;
        RECT 1539.130 2626.090 1540.310 2627.270 ;
        RECT 1540.730 2626.090 1541.910 2627.270 ;
        RECT 1539.130 2624.490 1540.310 2625.670 ;
        RECT 1540.730 2624.490 1541.910 2625.670 ;
        RECT 1539.130 2446.090 1540.310 2447.270 ;
        RECT 1540.730 2446.090 1541.910 2447.270 ;
        RECT 1539.130 2444.490 1540.310 2445.670 ;
        RECT 1540.730 2444.490 1541.910 2445.670 ;
        RECT 1539.130 2266.090 1540.310 2267.270 ;
        RECT 1540.730 2266.090 1541.910 2267.270 ;
        RECT 1539.130 2264.490 1540.310 2265.670 ;
        RECT 1540.730 2264.490 1541.910 2265.670 ;
        RECT 1539.130 2086.090 1540.310 2087.270 ;
        RECT 1540.730 2086.090 1541.910 2087.270 ;
        RECT 1539.130 2084.490 1540.310 2085.670 ;
        RECT 1540.730 2084.490 1541.910 2085.670 ;
        RECT 1539.130 1906.090 1540.310 1907.270 ;
        RECT 1540.730 1906.090 1541.910 1907.270 ;
        RECT 1539.130 1904.490 1540.310 1905.670 ;
        RECT 1540.730 1904.490 1541.910 1905.670 ;
        RECT 1539.130 1726.090 1540.310 1727.270 ;
        RECT 1540.730 1726.090 1541.910 1727.270 ;
        RECT 1539.130 1724.490 1540.310 1725.670 ;
        RECT 1540.730 1724.490 1541.910 1725.670 ;
        RECT 1539.130 1546.090 1540.310 1547.270 ;
        RECT 1540.730 1546.090 1541.910 1547.270 ;
        RECT 1539.130 1544.490 1540.310 1545.670 ;
        RECT 1540.730 1544.490 1541.910 1545.670 ;
        RECT 1539.130 1366.090 1540.310 1367.270 ;
        RECT 1540.730 1366.090 1541.910 1367.270 ;
        RECT 1539.130 1364.490 1540.310 1365.670 ;
        RECT 1540.730 1364.490 1541.910 1365.670 ;
        RECT 1539.130 1186.090 1540.310 1187.270 ;
        RECT 1540.730 1186.090 1541.910 1187.270 ;
        RECT 1539.130 1184.490 1540.310 1185.670 ;
        RECT 1540.730 1184.490 1541.910 1185.670 ;
        RECT 1539.130 1006.090 1540.310 1007.270 ;
        RECT 1540.730 1006.090 1541.910 1007.270 ;
        RECT 1539.130 1004.490 1540.310 1005.670 ;
        RECT 1540.730 1004.490 1541.910 1005.670 ;
        RECT 1539.130 826.090 1540.310 827.270 ;
        RECT 1540.730 826.090 1541.910 827.270 ;
        RECT 1539.130 824.490 1540.310 825.670 ;
        RECT 1540.730 824.490 1541.910 825.670 ;
        RECT 1539.130 646.090 1540.310 647.270 ;
        RECT 1540.730 646.090 1541.910 647.270 ;
        RECT 1539.130 644.490 1540.310 645.670 ;
        RECT 1540.730 644.490 1541.910 645.670 ;
        RECT 1539.130 466.090 1540.310 467.270 ;
        RECT 1540.730 466.090 1541.910 467.270 ;
        RECT 1539.130 464.490 1540.310 465.670 ;
        RECT 1540.730 464.490 1541.910 465.670 ;
        RECT 1539.130 286.090 1540.310 287.270 ;
        RECT 1540.730 286.090 1541.910 287.270 ;
        RECT 1539.130 284.490 1540.310 285.670 ;
        RECT 1540.730 284.490 1541.910 285.670 ;
        RECT 1539.130 106.090 1540.310 107.270 ;
        RECT 1540.730 106.090 1541.910 107.270 ;
        RECT 1539.130 104.490 1540.310 105.670 ;
        RECT 1540.730 104.490 1541.910 105.670 ;
        RECT 1539.130 -23.660 1540.310 -22.480 ;
        RECT 1540.730 -23.660 1541.910 -22.480 ;
        RECT 1539.130 -25.260 1540.310 -24.080 ;
        RECT 1540.730 -25.260 1541.910 -24.080 ;
        RECT 1719.130 3543.760 1720.310 3544.940 ;
        RECT 1720.730 3543.760 1721.910 3544.940 ;
        RECT 1719.130 3542.160 1720.310 3543.340 ;
        RECT 1720.730 3542.160 1721.910 3543.340 ;
        RECT 1719.130 3346.090 1720.310 3347.270 ;
        RECT 1720.730 3346.090 1721.910 3347.270 ;
        RECT 1719.130 3344.490 1720.310 3345.670 ;
        RECT 1720.730 3344.490 1721.910 3345.670 ;
        RECT 1719.130 3166.090 1720.310 3167.270 ;
        RECT 1720.730 3166.090 1721.910 3167.270 ;
        RECT 1719.130 3164.490 1720.310 3165.670 ;
        RECT 1720.730 3164.490 1721.910 3165.670 ;
        RECT 1719.130 2986.090 1720.310 2987.270 ;
        RECT 1720.730 2986.090 1721.910 2987.270 ;
        RECT 1719.130 2984.490 1720.310 2985.670 ;
        RECT 1720.730 2984.490 1721.910 2985.670 ;
        RECT 1719.130 2806.090 1720.310 2807.270 ;
        RECT 1720.730 2806.090 1721.910 2807.270 ;
        RECT 1719.130 2804.490 1720.310 2805.670 ;
        RECT 1720.730 2804.490 1721.910 2805.670 ;
        RECT 1719.130 2626.090 1720.310 2627.270 ;
        RECT 1720.730 2626.090 1721.910 2627.270 ;
        RECT 1719.130 2624.490 1720.310 2625.670 ;
        RECT 1720.730 2624.490 1721.910 2625.670 ;
        RECT 1719.130 2446.090 1720.310 2447.270 ;
        RECT 1720.730 2446.090 1721.910 2447.270 ;
        RECT 1719.130 2444.490 1720.310 2445.670 ;
        RECT 1720.730 2444.490 1721.910 2445.670 ;
        RECT 1719.130 2266.090 1720.310 2267.270 ;
        RECT 1720.730 2266.090 1721.910 2267.270 ;
        RECT 1719.130 2264.490 1720.310 2265.670 ;
        RECT 1720.730 2264.490 1721.910 2265.670 ;
        RECT 1719.130 2086.090 1720.310 2087.270 ;
        RECT 1720.730 2086.090 1721.910 2087.270 ;
        RECT 1719.130 2084.490 1720.310 2085.670 ;
        RECT 1720.730 2084.490 1721.910 2085.670 ;
        RECT 1719.130 1906.090 1720.310 1907.270 ;
        RECT 1720.730 1906.090 1721.910 1907.270 ;
        RECT 1719.130 1904.490 1720.310 1905.670 ;
        RECT 1720.730 1904.490 1721.910 1905.670 ;
        RECT 1719.130 1726.090 1720.310 1727.270 ;
        RECT 1720.730 1726.090 1721.910 1727.270 ;
        RECT 1719.130 1724.490 1720.310 1725.670 ;
        RECT 1720.730 1724.490 1721.910 1725.670 ;
        RECT 1719.130 1546.090 1720.310 1547.270 ;
        RECT 1720.730 1546.090 1721.910 1547.270 ;
        RECT 1719.130 1544.490 1720.310 1545.670 ;
        RECT 1720.730 1544.490 1721.910 1545.670 ;
        RECT 1719.130 1366.090 1720.310 1367.270 ;
        RECT 1720.730 1366.090 1721.910 1367.270 ;
        RECT 1719.130 1364.490 1720.310 1365.670 ;
        RECT 1720.730 1364.490 1721.910 1365.670 ;
        RECT 1719.130 1186.090 1720.310 1187.270 ;
        RECT 1720.730 1186.090 1721.910 1187.270 ;
        RECT 1719.130 1184.490 1720.310 1185.670 ;
        RECT 1720.730 1184.490 1721.910 1185.670 ;
        RECT 1719.130 1006.090 1720.310 1007.270 ;
        RECT 1720.730 1006.090 1721.910 1007.270 ;
        RECT 1719.130 1004.490 1720.310 1005.670 ;
        RECT 1720.730 1004.490 1721.910 1005.670 ;
        RECT 1719.130 826.090 1720.310 827.270 ;
        RECT 1720.730 826.090 1721.910 827.270 ;
        RECT 1719.130 824.490 1720.310 825.670 ;
        RECT 1720.730 824.490 1721.910 825.670 ;
        RECT 1719.130 646.090 1720.310 647.270 ;
        RECT 1720.730 646.090 1721.910 647.270 ;
        RECT 1719.130 644.490 1720.310 645.670 ;
        RECT 1720.730 644.490 1721.910 645.670 ;
        RECT 1719.130 466.090 1720.310 467.270 ;
        RECT 1720.730 466.090 1721.910 467.270 ;
        RECT 1719.130 464.490 1720.310 465.670 ;
        RECT 1720.730 464.490 1721.910 465.670 ;
        RECT 1719.130 286.090 1720.310 287.270 ;
        RECT 1720.730 286.090 1721.910 287.270 ;
        RECT 1719.130 284.490 1720.310 285.670 ;
        RECT 1720.730 284.490 1721.910 285.670 ;
        RECT 1719.130 106.090 1720.310 107.270 ;
        RECT 1720.730 106.090 1721.910 107.270 ;
        RECT 1719.130 104.490 1720.310 105.670 ;
        RECT 1720.730 104.490 1721.910 105.670 ;
        RECT 1719.130 -23.660 1720.310 -22.480 ;
        RECT 1720.730 -23.660 1721.910 -22.480 ;
        RECT 1719.130 -25.260 1720.310 -24.080 ;
        RECT 1720.730 -25.260 1721.910 -24.080 ;
        RECT 1899.130 3543.760 1900.310 3544.940 ;
        RECT 1900.730 3543.760 1901.910 3544.940 ;
        RECT 1899.130 3542.160 1900.310 3543.340 ;
        RECT 1900.730 3542.160 1901.910 3543.340 ;
        RECT 1899.130 3346.090 1900.310 3347.270 ;
        RECT 1900.730 3346.090 1901.910 3347.270 ;
        RECT 1899.130 3344.490 1900.310 3345.670 ;
        RECT 1900.730 3344.490 1901.910 3345.670 ;
        RECT 1899.130 3166.090 1900.310 3167.270 ;
        RECT 1900.730 3166.090 1901.910 3167.270 ;
        RECT 1899.130 3164.490 1900.310 3165.670 ;
        RECT 1900.730 3164.490 1901.910 3165.670 ;
        RECT 1899.130 2986.090 1900.310 2987.270 ;
        RECT 1900.730 2986.090 1901.910 2987.270 ;
        RECT 1899.130 2984.490 1900.310 2985.670 ;
        RECT 1900.730 2984.490 1901.910 2985.670 ;
        RECT 1899.130 2806.090 1900.310 2807.270 ;
        RECT 1900.730 2806.090 1901.910 2807.270 ;
        RECT 1899.130 2804.490 1900.310 2805.670 ;
        RECT 1900.730 2804.490 1901.910 2805.670 ;
        RECT 1899.130 2626.090 1900.310 2627.270 ;
        RECT 1900.730 2626.090 1901.910 2627.270 ;
        RECT 1899.130 2624.490 1900.310 2625.670 ;
        RECT 1900.730 2624.490 1901.910 2625.670 ;
        RECT 1899.130 2446.090 1900.310 2447.270 ;
        RECT 1900.730 2446.090 1901.910 2447.270 ;
        RECT 1899.130 2444.490 1900.310 2445.670 ;
        RECT 1900.730 2444.490 1901.910 2445.670 ;
        RECT 1899.130 2266.090 1900.310 2267.270 ;
        RECT 1900.730 2266.090 1901.910 2267.270 ;
        RECT 1899.130 2264.490 1900.310 2265.670 ;
        RECT 1900.730 2264.490 1901.910 2265.670 ;
        RECT 1899.130 2086.090 1900.310 2087.270 ;
        RECT 1900.730 2086.090 1901.910 2087.270 ;
        RECT 1899.130 2084.490 1900.310 2085.670 ;
        RECT 1900.730 2084.490 1901.910 2085.670 ;
        RECT 1899.130 1906.090 1900.310 1907.270 ;
        RECT 1900.730 1906.090 1901.910 1907.270 ;
        RECT 1899.130 1904.490 1900.310 1905.670 ;
        RECT 1900.730 1904.490 1901.910 1905.670 ;
        RECT 1899.130 1726.090 1900.310 1727.270 ;
        RECT 1900.730 1726.090 1901.910 1727.270 ;
        RECT 1899.130 1724.490 1900.310 1725.670 ;
        RECT 1900.730 1724.490 1901.910 1725.670 ;
        RECT 1899.130 1546.090 1900.310 1547.270 ;
        RECT 1900.730 1546.090 1901.910 1547.270 ;
        RECT 1899.130 1544.490 1900.310 1545.670 ;
        RECT 1900.730 1544.490 1901.910 1545.670 ;
        RECT 1899.130 1366.090 1900.310 1367.270 ;
        RECT 1900.730 1366.090 1901.910 1367.270 ;
        RECT 1899.130 1364.490 1900.310 1365.670 ;
        RECT 1900.730 1364.490 1901.910 1365.670 ;
        RECT 1899.130 1186.090 1900.310 1187.270 ;
        RECT 1900.730 1186.090 1901.910 1187.270 ;
        RECT 1899.130 1184.490 1900.310 1185.670 ;
        RECT 1900.730 1184.490 1901.910 1185.670 ;
        RECT 1899.130 1006.090 1900.310 1007.270 ;
        RECT 1900.730 1006.090 1901.910 1007.270 ;
        RECT 1899.130 1004.490 1900.310 1005.670 ;
        RECT 1900.730 1004.490 1901.910 1005.670 ;
        RECT 1899.130 826.090 1900.310 827.270 ;
        RECT 1900.730 826.090 1901.910 827.270 ;
        RECT 1899.130 824.490 1900.310 825.670 ;
        RECT 1900.730 824.490 1901.910 825.670 ;
        RECT 1899.130 646.090 1900.310 647.270 ;
        RECT 1900.730 646.090 1901.910 647.270 ;
        RECT 1899.130 644.490 1900.310 645.670 ;
        RECT 1900.730 644.490 1901.910 645.670 ;
        RECT 1899.130 466.090 1900.310 467.270 ;
        RECT 1900.730 466.090 1901.910 467.270 ;
        RECT 1899.130 464.490 1900.310 465.670 ;
        RECT 1900.730 464.490 1901.910 465.670 ;
        RECT 1899.130 286.090 1900.310 287.270 ;
        RECT 1900.730 286.090 1901.910 287.270 ;
        RECT 1899.130 284.490 1900.310 285.670 ;
        RECT 1900.730 284.490 1901.910 285.670 ;
        RECT 1899.130 106.090 1900.310 107.270 ;
        RECT 1900.730 106.090 1901.910 107.270 ;
        RECT 1899.130 104.490 1900.310 105.670 ;
        RECT 1900.730 104.490 1901.910 105.670 ;
        RECT 1899.130 -23.660 1900.310 -22.480 ;
        RECT 1900.730 -23.660 1901.910 -22.480 ;
        RECT 1899.130 -25.260 1900.310 -24.080 ;
        RECT 1900.730 -25.260 1901.910 -24.080 ;
        RECT 2079.130 3543.760 2080.310 3544.940 ;
        RECT 2080.730 3543.760 2081.910 3544.940 ;
        RECT 2079.130 3542.160 2080.310 3543.340 ;
        RECT 2080.730 3542.160 2081.910 3543.340 ;
        RECT 2079.130 3346.090 2080.310 3347.270 ;
        RECT 2080.730 3346.090 2081.910 3347.270 ;
        RECT 2079.130 3344.490 2080.310 3345.670 ;
        RECT 2080.730 3344.490 2081.910 3345.670 ;
        RECT 2079.130 3166.090 2080.310 3167.270 ;
        RECT 2080.730 3166.090 2081.910 3167.270 ;
        RECT 2079.130 3164.490 2080.310 3165.670 ;
        RECT 2080.730 3164.490 2081.910 3165.670 ;
        RECT 2079.130 2986.090 2080.310 2987.270 ;
        RECT 2080.730 2986.090 2081.910 2987.270 ;
        RECT 2079.130 2984.490 2080.310 2985.670 ;
        RECT 2080.730 2984.490 2081.910 2985.670 ;
        RECT 2079.130 2806.090 2080.310 2807.270 ;
        RECT 2080.730 2806.090 2081.910 2807.270 ;
        RECT 2079.130 2804.490 2080.310 2805.670 ;
        RECT 2080.730 2804.490 2081.910 2805.670 ;
        RECT 2079.130 2626.090 2080.310 2627.270 ;
        RECT 2080.730 2626.090 2081.910 2627.270 ;
        RECT 2079.130 2624.490 2080.310 2625.670 ;
        RECT 2080.730 2624.490 2081.910 2625.670 ;
        RECT 2079.130 2446.090 2080.310 2447.270 ;
        RECT 2080.730 2446.090 2081.910 2447.270 ;
        RECT 2079.130 2444.490 2080.310 2445.670 ;
        RECT 2080.730 2444.490 2081.910 2445.670 ;
        RECT 2079.130 2266.090 2080.310 2267.270 ;
        RECT 2080.730 2266.090 2081.910 2267.270 ;
        RECT 2079.130 2264.490 2080.310 2265.670 ;
        RECT 2080.730 2264.490 2081.910 2265.670 ;
        RECT 2079.130 2086.090 2080.310 2087.270 ;
        RECT 2080.730 2086.090 2081.910 2087.270 ;
        RECT 2079.130 2084.490 2080.310 2085.670 ;
        RECT 2080.730 2084.490 2081.910 2085.670 ;
        RECT 2079.130 1906.090 2080.310 1907.270 ;
        RECT 2080.730 1906.090 2081.910 1907.270 ;
        RECT 2079.130 1904.490 2080.310 1905.670 ;
        RECT 2080.730 1904.490 2081.910 1905.670 ;
        RECT 2079.130 1726.090 2080.310 1727.270 ;
        RECT 2080.730 1726.090 2081.910 1727.270 ;
        RECT 2079.130 1724.490 2080.310 1725.670 ;
        RECT 2080.730 1724.490 2081.910 1725.670 ;
        RECT 2079.130 1546.090 2080.310 1547.270 ;
        RECT 2080.730 1546.090 2081.910 1547.270 ;
        RECT 2079.130 1544.490 2080.310 1545.670 ;
        RECT 2080.730 1544.490 2081.910 1545.670 ;
        RECT 2079.130 1366.090 2080.310 1367.270 ;
        RECT 2080.730 1366.090 2081.910 1367.270 ;
        RECT 2079.130 1364.490 2080.310 1365.670 ;
        RECT 2080.730 1364.490 2081.910 1365.670 ;
        RECT 2079.130 1186.090 2080.310 1187.270 ;
        RECT 2080.730 1186.090 2081.910 1187.270 ;
        RECT 2079.130 1184.490 2080.310 1185.670 ;
        RECT 2080.730 1184.490 2081.910 1185.670 ;
        RECT 2079.130 1006.090 2080.310 1007.270 ;
        RECT 2080.730 1006.090 2081.910 1007.270 ;
        RECT 2079.130 1004.490 2080.310 1005.670 ;
        RECT 2080.730 1004.490 2081.910 1005.670 ;
        RECT 2079.130 826.090 2080.310 827.270 ;
        RECT 2080.730 826.090 2081.910 827.270 ;
        RECT 2079.130 824.490 2080.310 825.670 ;
        RECT 2080.730 824.490 2081.910 825.670 ;
        RECT 2079.130 646.090 2080.310 647.270 ;
        RECT 2080.730 646.090 2081.910 647.270 ;
        RECT 2079.130 644.490 2080.310 645.670 ;
        RECT 2080.730 644.490 2081.910 645.670 ;
        RECT 2079.130 466.090 2080.310 467.270 ;
        RECT 2080.730 466.090 2081.910 467.270 ;
        RECT 2079.130 464.490 2080.310 465.670 ;
        RECT 2080.730 464.490 2081.910 465.670 ;
        RECT 2079.130 286.090 2080.310 287.270 ;
        RECT 2080.730 286.090 2081.910 287.270 ;
        RECT 2079.130 284.490 2080.310 285.670 ;
        RECT 2080.730 284.490 2081.910 285.670 ;
        RECT 2079.130 106.090 2080.310 107.270 ;
        RECT 2080.730 106.090 2081.910 107.270 ;
        RECT 2079.130 104.490 2080.310 105.670 ;
        RECT 2080.730 104.490 2081.910 105.670 ;
        RECT 2079.130 -23.660 2080.310 -22.480 ;
        RECT 2080.730 -23.660 2081.910 -22.480 ;
        RECT 2079.130 -25.260 2080.310 -24.080 ;
        RECT 2080.730 -25.260 2081.910 -24.080 ;
        RECT 2259.130 3543.760 2260.310 3544.940 ;
        RECT 2260.730 3543.760 2261.910 3544.940 ;
        RECT 2259.130 3542.160 2260.310 3543.340 ;
        RECT 2260.730 3542.160 2261.910 3543.340 ;
        RECT 2259.130 3346.090 2260.310 3347.270 ;
        RECT 2260.730 3346.090 2261.910 3347.270 ;
        RECT 2259.130 3344.490 2260.310 3345.670 ;
        RECT 2260.730 3344.490 2261.910 3345.670 ;
        RECT 2259.130 3166.090 2260.310 3167.270 ;
        RECT 2260.730 3166.090 2261.910 3167.270 ;
        RECT 2259.130 3164.490 2260.310 3165.670 ;
        RECT 2260.730 3164.490 2261.910 3165.670 ;
        RECT 2259.130 2986.090 2260.310 2987.270 ;
        RECT 2260.730 2986.090 2261.910 2987.270 ;
        RECT 2259.130 2984.490 2260.310 2985.670 ;
        RECT 2260.730 2984.490 2261.910 2985.670 ;
        RECT 2259.130 2806.090 2260.310 2807.270 ;
        RECT 2260.730 2806.090 2261.910 2807.270 ;
        RECT 2259.130 2804.490 2260.310 2805.670 ;
        RECT 2260.730 2804.490 2261.910 2805.670 ;
        RECT 2259.130 2626.090 2260.310 2627.270 ;
        RECT 2260.730 2626.090 2261.910 2627.270 ;
        RECT 2259.130 2624.490 2260.310 2625.670 ;
        RECT 2260.730 2624.490 2261.910 2625.670 ;
        RECT 2259.130 2446.090 2260.310 2447.270 ;
        RECT 2260.730 2446.090 2261.910 2447.270 ;
        RECT 2259.130 2444.490 2260.310 2445.670 ;
        RECT 2260.730 2444.490 2261.910 2445.670 ;
        RECT 2259.130 2266.090 2260.310 2267.270 ;
        RECT 2260.730 2266.090 2261.910 2267.270 ;
        RECT 2259.130 2264.490 2260.310 2265.670 ;
        RECT 2260.730 2264.490 2261.910 2265.670 ;
        RECT 2259.130 2086.090 2260.310 2087.270 ;
        RECT 2260.730 2086.090 2261.910 2087.270 ;
        RECT 2259.130 2084.490 2260.310 2085.670 ;
        RECT 2260.730 2084.490 2261.910 2085.670 ;
        RECT 2259.130 1906.090 2260.310 1907.270 ;
        RECT 2260.730 1906.090 2261.910 1907.270 ;
        RECT 2259.130 1904.490 2260.310 1905.670 ;
        RECT 2260.730 1904.490 2261.910 1905.670 ;
        RECT 2259.130 1726.090 2260.310 1727.270 ;
        RECT 2260.730 1726.090 2261.910 1727.270 ;
        RECT 2259.130 1724.490 2260.310 1725.670 ;
        RECT 2260.730 1724.490 2261.910 1725.670 ;
        RECT 2259.130 1546.090 2260.310 1547.270 ;
        RECT 2260.730 1546.090 2261.910 1547.270 ;
        RECT 2259.130 1544.490 2260.310 1545.670 ;
        RECT 2260.730 1544.490 2261.910 1545.670 ;
        RECT 2259.130 1366.090 2260.310 1367.270 ;
        RECT 2260.730 1366.090 2261.910 1367.270 ;
        RECT 2259.130 1364.490 2260.310 1365.670 ;
        RECT 2260.730 1364.490 2261.910 1365.670 ;
        RECT 2259.130 1186.090 2260.310 1187.270 ;
        RECT 2260.730 1186.090 2261.910 1187.270 ;
        RECT 2259.130 1184.490 2260.310 1185.670 ;
        RECT 2260.730 1184.490 2261.910 1185.670 ;
        RECT 2259.130 1006.090 2260.310 1007.270 ;
        RECT 2260.730 1006.090 2261.910 1007.270 ;
        RECT 2259.130 1004.490 2260.310 1005.670 ;
        RECT 2260.730 1004.490 2261.910 1005.670 ;
        RECT 2259.130 826.090 2260.310 827.270 ;
        RECT 2260.730 826.090 2261.910 827.270 ;
        RECT 2259.130 824.490 2260.310 825.670 ;
        RECT 2260.730 824.490 2261.910 825.670 ;
        RECT 2259.130 646.090 2260.310 647.270 ;
        RECT 2260.730 646.090 2261.910 647.270 ;
        RECT 2259.130 644.490 2260.310 645.670 ;
        RECT 2260.730 644.490 2261.910 645.670 ;
        RECT 2259.130 466.090 2260.310 467.270 ;
        RECT 2260.730 466.090 2261.910 467.270 ;
        RECT 2259.130 464.490 2260.310 465.670 ;
        RECT 2260.730 464.490 2261.910 465.670 ;
        RECT 2259.130 286.090 2260.310 287.270 ;
        RECT 2260.730 286.090 2261.910 287.270 ;
        RECT 2259.130 284.490 2260.310 285.670 ;
        RECT 2260.730 284.490 2261.910 285.670 ;
        RECT 2259.130 106.090 2260.310 107.270 ;
        RECT 2260.730 106.090 2261.910 107.270 ;
        RECT 2259.130 104.490 2260.310 105.670 ;
        RECT 2260.730 104.490 2261.910 105.670 ;
        RECT 2259.130 -23.660 2260.310 -22.480 ;
        RECT 2260.730 -23.660 2261.910 -22.480 ;
        RECT 2259.130 -25.260 2260.310 -24.080 ;
        RECT 2260.730 -25.260 2261.910 -24.080 ;
        RECT 2439.130 3543.760 2440.310 3544.940 ;
        RECT 2440.730 3543.760 2441.910 3544.940 ;
        RECT 2439.130 3542.160 2440.310 3543.340 ;
        RECT 2440.730 3542.160 2441.910 3543.340 ;
        RECT 2439.130 3346.090 2440.310 3347.270 ;
        RECT 2440.730 3346.090 2441.910 3347.270 ;
        RECT 2439.130 3344.490 2440.310 3345.670 ;
        RECT 2440.730 3344.490 2441.910 3345.670 ;
        RECT 2439.130 3166.090 2440.310 3167.270 ;
        RECT 2440.730 3166.090 2441.910 3167.270 ;
        RECT 2439.130 3164.490 2440.310 3165.670 ;
        RECT 2440.730 3164.490 2441.910 3165.670 ;
        RECT 2439.130 2986.090 2440.310 2987.270 ;
        RECT 2440.730 2986.090 2441.910 2987.270 ;
        RECT 2439.130 2984.490 2440.310 2985.670 ;
        RECT 2440.730 2984.490 2441.910 2985.670 ;
        RECT 2439.130 2806.090 2440.310 2807.270 ;
        RECT 2440.730 2806.090 2441.910 2807.270 ;
        RECT 2439.130 2804.490 2440.310 2805.670 ;
        RECT 2440.730 2804.490 2441.910 2805.670 ;
        RECT 2439.130 2626.090 2440.310 2627.270 ;
        RECT 2440.730 2626.090 2441.910 2627.270 ;
        RECT 2439.130 2624.490 2440.310 2625.670 ;
        RECT 2440.730 2624.490 2441.910 2625.670 ;
        RECT 2439.130 2446.090 2440.310 2447.270 ;
        RECT 2440.730 2446.090 2441.910 2447.270 ;
        RECT 2439.130 2444.490 2440.310 2445.670 ;
        RECT 2440.730 2444.490 2441.910 2445.670 ;
        RECT 2439.130 2266.090 2440.310 2267.270 ;
        RECT 2440.730 2266.090 2441.910 2267.270 ;
        RECT 2439.130 2264.490 2440.310 2265.670 ;
        RECT 2440.730 2264.490 2441.910 2265.670 ;
        RECT 2439.130 2086.090 2440.310 2087.270 ;
        RECT 2440.730 2086.090 2441.910 2087.270 ;
        RECT 2439.130 2084.490 2440.310 2085.670 ;
        RECT 2440.730 2084.490 2441.910 2085.670 ;
        RECT 2439.130 1906.090 2440.310 1907.270 ;
        RECT 2440.730 1906.090 2441.910 1907.270 ;
        RECT 2439.130 1904.490 2440.310 1905.670 ;
        RECT 2440.730 1904.490 2441.910 1905.670 ;
        RECT 2439.130 1726.090 2440.310 1727.270 ;
        RECT 2440.730 1726.090 2441.910 1727.270 ;
        RECT 2439.130 1724.490 2440.310 1725.670 ;
        RECT 2440.730 1724.490 2441.910 1725.670 ;
        RECT 2439.130 1546.090 2440.310 1547.270 ;
        RECT 2440.730 1546.090 2441.910 1547.270 ;
        RECT 2439.130 1544.490 2440.310 1545.670 ;
        RECT 2440.730 1544.490 2441.910 1545.670 ;
        RECT 2439.130 1366.090 2440.310 1367.270 ;
        RECT 2440.730 1366.090 2441.910 1367.270 ;
        RECT 2439.130 1364.490 2440.310 1365.670 ;
        RECT 2440.730 1364.490 2441.910 1365.670 ;
        RECT 2439.130 1186.090 2440.310 1187.270 ;
        RECT 2440.730 1186.090 2441.910 1187.270 ;
        RECT 2439.130 1184.490 2440.310 1185.670 ;
        RECT 2440.730 1184.490 2441.910 1185.670 ;
        RECT 2439.130 1006.090 2440.310 1007.270 ;
        RECT 2440.730 1006.090 2441.910 1007.270 ;
        RECT 2439.130 1004.490 2440.310 1005.670 ;
        RECT 2440.730 1004.490 2441.910 1005.670 ;
        RECT 2439.130 826.090 2440.310 827.270 ;
        RECT 2440.730 826.090 2441.910 827.270 ;
        RECT 2439.130 824.490 2440.310 825.670 ;
        RECT 2440.730 824.490 2441.910 825.670 ;
        RECT 2439.130 646.090 2440.310 647.270 ;
        RECT 2440.730 646.090 2441.910 647.270 ;
        RECT 2439.130 644.490 2440.310 645.670 ;
        RECT 2440.730 644.490 2441.910 645.670 ;
        RECT 2439.130 466.090 2440.310 467.270 ;
        RECT 2440.730 466.090 2441.910 467.270 ;
        RECT 2439.130 464.490 2440.310 465.670 ;
        RECT 2440.730 464.490 2441.910 465.670 ;
        RECT 2439.130 286.090 2440.310 287.270 ;
        RECT 2440.730 286.090 2441.910 287.270 ;
        RECT 2439.130 284.490 2440.310 285.670 ;
        RECT 2440.730 284.490 2441.910 285.670 ;
        RECT 2439.130 106.090 2440.310 107.270 ;
        RECT 2440.730 106.090 2441.910 107.270 ;
        RECT 2439.130 104.490 2440.310 105.670 ;
        RECT 2440.730 104.490 2441.910 105.670 ;
        RECT 2439.130 -23.660 2440.310 -22.480 ;
        RECT 2440.730 -23.660 2441.910 -22.480 ;
        RECT 2439.130 -25.260 2440.310 -24.080 ;
        RECT 2440.730 -25.260 2441.910 -24.080 ;
        RECT 2619.130 3543.760 2620.310 3544.940 ;
        RECT 2620.730 3543.760 2621.910 3544.940 ;
        RECT 2619.130 3542.160 2620.310 3543.340 ;
        RECT 2620.730 3542.160 2621.910 3543.340 ;
        RECT 2619.130 3346.090 2620.310 3347.270 ;
        RECT 2620.730 3346.090 2621.910 3347.270 ;
        RECT 2619.130 3344.490 2620.310 3345.670 ;
        RECT 2620.730 3344.490 2621.910 3345.670 ;
        RECT 2619.130 3166.090 2620.310 3167.270 ;
        RECT 2620.730 3166.090 2621.910 3167.270 ;
        RECT 2619.130 3164.490 2620.310 3165.670 ;
        RECT 2620.730 3164.490 2621.910 3165.670 ;
        RECT 2619.130 2986.090 2620.310 2987.270 ;
        RECT 2620.730 2986.090 2621.910 2987.270 ;
        RECT 2619.130 2984.490 2620.310 2985.670 ;
        RECT 2620.730 2984.490 2621.910 2985.670 ;
        RECT 2619.130 2806.090 2620.310 2807.270 ;
        RECT 2620.730 2806.090 2621.910 2807.270 ;
        RECT 2619.130 2804.490 2620.310 2805.670 ;
        RECT 2620.730 2804.490 2621.910 2805.670 ;
        RECT 2619.130 2626.090 2620.310 2627.270 ;
        RECT 2620.730 2626.090 2621.910 2627.270 ;
        RECT 2619.130 2624.490 2620.310 2625.670 ;
        RECT 2620.730 2624.490 2621.910 2625.670 ;
        RECT 2619.130 2446.090 2620.310 2447.270 ;
        RECT 2620.730 2446.090 2621.910 2447.270 ;
        RECT 2619.130 2444.490 2620.310 2445.670 ;
        RECT 2620.730 2444.490 2621.910 2445.670 ;
        RECT 2619.130 2266.090 2620.310 2267.270 ;
        RECT 2620.730 2266.090 2621.910 2267.270 ;
        RECT 2619.130 2264.490 2620.310 2265.670 ;
        RECT 2620.730 2264.490 2621.910 2265.670 ;
        RECT 2619.130 2086.090 2620.310 2087.270 ;
        RECT 2620.730 2086.090 2621.910 2087.270 ;
        RECT 2619.130 2084.490 2620.310 2085.670 ;
        RECT 2620.730 2084.490 2621.910 2085.670 ;
        RECT 2619.130 1906.090 2620.310 1907.270 ;
        RECT 2620.730 1906.090 2621.910 1907.270 ;
        RECT 2619.130 1904.490 2620.310 1905.670 ;
        RECT 2620.730 1904.490 2621.910 1905.670 ;
        RECT 2619.130 1726.090 2620.310 1727.270 ;
        RECT 2620.730 1726.090 2621.910 1727.270 ;
        RECT 2619.130 1724.490 2620.310 1725.670 ;
        RECT 2620.730 1724.490 2621.910 1725.670 ;
        RECT 2619.130 1546.090 2620.310 1547.270 ;
        RECT 2620.730 1546.090 2621.910 1547.270 ;
        RECT 2619.130 1544.490 2620.310 1545.670 ;
        RECT 2620.730 1544.490 2621.910 1545.670 ;
        RECT 2619.130 1366.090 2620.310 1367.270 ;
        RECT 2620.730 1366.090 2621.910 1367.270 ;
        RECT 2619.130 1364.490 2620.310 1365.670 ;
        RECT 2620.730 1364.490 2621.910 1365.670 ;
        RECT 2619.130 1186.090 2620.310 1187.270 ;
        RECT 2620.730 1186.090 2621.910 1187.270 ;
        RECT 2619.130 1184.490 2620.310 1185.670 ;
        RECT 2620.730 1184.490 2621.910 1185.670 ;
        RECT 2619.130 1006.090 2620.310 1007.270 ;
        RECT 2620.730 1006.090 2621.910 1007.270 ;
        RECT 2619.130 1004.490 2620.310 1005.670 ;
        RECT 2620.730 1004.490 2621.910 1005.670 ;
        RECT 2619.130 826.090 2620.310 827.270 ;
        RECT 2620.730 826.090 2621.910 827.270 ;
        RECT 2619.130 824.490 2620.310 825.670 ;
        RECT 2620.730 824.490 2621.910 825.670 ;
        RECT 2619.130 646.090 2620.310 647.270 ;
        RECT 2620.730 646.090 2621.910 647.270 ;
        RECT 2619.130 644.490 2620.310 645.670 ;
        RECT 2620.730 644.490 2621.910 645.670 ;
        RECT 2619.130 466.090 2620.310 467.270 ;
        RECT 2620.730 466.090 2621.910 467.270 ;
        RECT 2619.130 464.490 2620.310 465.670 ;
        RECT 2620.730 464.490 2621.910 465.670 ;
        RECT 2619.130 286.090 2620.310 287.270 ;
        RECT 2620.730 286.090 2621.910 287.270 ;
        RECT 2619.130 284.490 2620.310 285.670 ;
        RECT 2620.730 284.490 2621.910 285.670 ;
        RECT 2619.130 106.090 2620.310 107.270 ;
        RECT 2620.730 106.090 2621.910 107.270 ;
        RECT 2619.130 104.490 2620.310 105.670 ;
        RECT 2620.730 104.490 2621.910 105.670 ;
        RECT 2619.130 -23.660 2620.310 -22.480 ;
        RECT 2620.730 -23.660 2621.910 -22.480 ;
        RECT 2619.130 -25.260 2620.310 -24.080 ;
        RECT 2620.730 -25.260 2621.910 -24.080 ;
        RECT 2799.130 3543.760 2800.310 3544.940 ;
        RECT 2800.730 3543.760 2801.910 3544.940 ;
        RECT 2799.130 3542.160 2800.310 3543.340 ;
        RECT 2800.730 3542.160 2801.910 3543.340 ;
        RECT 2799.130 3346.090 2800.310 3347.270 ;
        RECT 2800.730 3346.090 2801.910 3347.270 ;
        RECT 2799.130 3344.490 2800.310 3345.670 ;
        RECT 2800.730 3344.490 2801.910 3345.670 ;
        RECT 2799.130 3166.090 2800.310 3167.270 ;
        RECT 2800.730 3166.090 2801.910 3167.270 ;
        RECT 2799.130 3164.490 2800.310 3165.670 ;
        RECT 2800.730 3164.490 2801.910 3165.670 ;
        RECT 2799.130 2986.090 2800.310 2987.270 ;
        RECT 2800.730 2986.090 2801.910 2987.270 ;
        RECT 2799.130 2984.490 2800.310 2985.670 ;
        RECT 2800.730 2984.490 2801.910 2985.670 ;
        RECT 2799.130 2806.090 2800.310 2807.270 ;
        RECT 2800.730 2806.090 2801.910 2807.270 ;
        RECT 2799.130 2804.490 2800.310 2805.670 ;
        RECT 2800.730 2804.490 2801.910 2805.670 ;
        RECT 2799.130 2626.090 2800.310 2627.270 ;
        RECT 2800.730 2626.090 2801.910 2627.270 ;
        RECT 2799.130 2624.490 2800.310 2625.670 ;
        RECT 2800.730 2624.490 2801.910 2625.670 ;
        RECT 2799.130 2446.090 2800.310 2447.270 ;
        RECT 2800.730 2446.090 2801.910 2447.270 ;
        RECT 2799.130 2444.490 2800.310 2445.670 ;
        RECT 2800.730 2444.490 2801.910 2445.670 ;
        RECT 2799.130 2266.090 2800.310 2267.270 ;
        RECT 2800.730 2266.090 2801.910 2267.270 ;
        RECT 2799.130 2264.490 2800.310 2265.670 ;
        RECT 2800.730 2264.490 2801.910 2265.670 ;
        RECT 2799.130 2086.090 2800.310 2087.270 ;
        RECT 2800.730 2086.090 2801.910 2087.270 ;
        RECT 2799.130 2084.490 2800.310 2085.670 ;
        RECT 2800.730 2084.490 2801.910 2085.670 ;
        RECT 2799.130 1906.090 2800.310 1907.270 ;
        RECT 2800.730 1906.090 2801.910 1907.270 ;
        RECT 2799.130 1904.490 2800.310 1905.670 ;
        RECT 2800.730 1904.490 2801.910 1905.670 ;
        RECT 2799.130 1726.090 2800.310 1727.270 ;
        RECT 2800.730 1726.090 2801.910 1727.270 ;
        RECT 2799.130 1724.490 2800.310 1725.670 ;
        RECT 2800.730 1724.490 2801.910 1725.670 ;
        RECT 2799.130 1546.090 2800.310 1547.270 ;
        RECT 2800.730 1546.090 2801.910 1547.270 ;
        RECT 2799.130 1544.490 2800.310 1545.670 ;
        RECT 2800.730 1544.490 2801.910 1545.670 ;
        RECT 2799.130 1366.090 2800.310 1367.270 ;
        RECT 2800.730 1366.090 2801.910 1367.270 ;
        RECT 2799.130 1364.490 2800.310 1365.670 ;
        RECT 2800.730 1364.490 2801.910 1365.670 ;
        RECT 2799.130 1186.090 2800.310 1187.270 ;
        RECT 2800.730 1186.090 2801.910 1187.270 ;
        RECT 2799.130 1184.490 2800.310 1185.670 ;
        RECT 2800.730 1184.490 2801.910 1185.670 ;
        RECT 2799.130 1006.090 2800.310 1007.270 ;
        RECT 2800.730 1006.090 2801.910 1007.270 ;
        RECT 2799.130 1004.490 2800.310 1005.670 ;
        RECT 2800.730 1004.490 2801.910 1005.670 ;
        RECT 2799.130 826.090 2800.310 827.270 ;
        RECT 2800.730 826.090 2801.910 827.270 ;
        RECT 2799.130 824.490 2800.310 825.670 ;
        RECT 2800.730 824.490 2801.910 825.670 ;
        RECT 2799.130 646.090 2800.310 647.270 ;
        RECT 2800.730 646.090 2801.910 647.270 ;
        RECT 2799.130 644.490 2800.310 645.670 ;
        RECT 2800.730 644.490 2801.910 645.670 ;
        RECT 2799.130 466.090 2800.310 467.270 ;
        RECT 2800.730 466.090 2801.910 467.270 ;
        RECT 2799.130 464.490 2800.310 465.670 ;
        RECT 2800.730 464.490 2801.910 465.670 ;
        RECT 2799.130 286.090 2800.310 287.270 ;
        RECT 2800.730 286.090 2801.910 287.270 ;
        RECT 2799.130 284.490 2800.310 285.670 ;
        RECT 2800.730 284.490 2801.910 285.670 ;
        RECT 2799.130 106.090 2800.310 107.270 ;
        RECT 2800.730 106.090 2801.910 107.270 ;
        RECT 2799.130 104.490 2800.310 105.670 ;
        RECT 2800.730 104.490 2801.910 105.670 ;
        RECT 2799.130 -23.660 2800.310 -22.480 ;
        RECT 2800.730 -23.660 2801.910 -22.480 ;
        RECT 2799.130 -25.260 2800.310 -24.080 ;
        RECT 2800.730 -25.260 2801.910 -24.080 ;
        RECT 2947.460 3543.760 2948.640 3544.940 ;
        RECT 2949.060 3543.760 2950.240 3544.940 ;
        RECT 2947.460 3542.160 2948.640 3543.340 ;
        RECT 2949.060 3542.160 2950.240 3543.340 ;
        RECT 2947.460 3346.090 2948.640 3347.270 ;
        RECT 2949.060 3346.090 2950.240 3347.270 ;
        RECT 2947.460 3344.490 2948.640 3345.670 ;
        RECT 2949.060 3344.490 2950.240 3345.670 ;
        RECT 2947.460 3166.090 2948.640 3167.270 ;
        RECT 2949.060 3166.090 2950.240 3167.270 ;
        RECT 2947.460 3164.490 2948.640 3165.670 ;
        RECT 2949.060 3164.490 2950.240 3165.670 ;
        RECT 2947.460 2986.090 2948.640 2987.270 ;
        RECT 2949.060 2986.090 2950.240 2987.270 ;
        RECT 2947.460 2984.490 2948.640 2985.670 ;
        RECT 2949.060 2984.490 2950.240 2985.670 ;
        RECT 2947.460 2806.090 2948.640 2807.270 ;
        RECT 2949.060 2806.090 2950.240 2807.270 ;
        RECT 2947.460 2804.490 2948.640 2805.670 ;
        RECT 2949.060 2804.490 2950.240 2805.670 ;
        RECT 2947.460 2626.090 2948.640 2627.270 ;
        RECT 2949.060 2626.090 2950.240 2627.270 ;
        RECT 2947.460 2624.490 2948.640 2625.670 ;
        RECT 2949.060 2624.490 2950.240 2625.670 ;
        RECT 2947.460 2446.090 2948.640 2447.270 ;
        RECT 2949.060 2446.090 2950.240 2447.270 ;
        RECT 2947.460 2444.490 2948.640 2445.670 ;
        RECT 2949.060 2444.490 2950.240 2445.670 ;
        RECT 2947.460 2266.090 2948.640 2267.270 ;
        RECT 2949.060 2266.090 2950.240 2267.270 ;
        RECT 2947.460 2264.490 2948.640 2265.670 ;
        RECT 2949.060 2264.490 2950.240 2265.670 ;
        RECT 2947.460 2086.090 2948.640 2087.270 ;
        RECT 2949.060 2086.090 2950.240 2087.270 ;
        RECT 2947.460 2084.490 2948.640 2085.670 ;
        RECT 2949.060 2084.490 2950.240 2085.670 ;
        RECT 2947.460 1906.090 2948.640 1907.270 ;
        RECT 2949.060 1906.090 2950.240 1907.270 ;
        RECT 2947.460 1904.490 2948.640 1905.670 ;
        RECT 2949.060 1904.490 2950.240 1905.670 ;
        RECT 2947.460 1726.090 2948.640 1727.270 ;
        RECT 2949.060 1726.090 2950.240 1727.270 ;
        RECT 2947.460 1724.490 2948.640 1725.670 ;
        RECT 2949.060 1724.490 2950.240 1725.670 ;
        RECT 2947.460 1546.090 2948.640 1547.270 ;
        RECT 2949.060 1546.090 2950.240 1547.270 ;
        RECT 2947.460 1544.490 2948.640 1545.670 ;
        RECT 2949.060 1544.490 2950.240 1545.670 ;
        RECT 2947.460 1366.090 2948.640 1367.270 ;
        RECT 2949.060 1366.090 2950.240 1367.270 ;
        RECT 2947.460 1364.490 2948.640 1365.670 ;
        RECT 2949.060 1364.490 2950.240 1365.670 ;
        RECT 2947.460 1186.090 2948.640 1187.270 ;
        RECT 2949.060 1186.090 2950.240 1187.270 ;
        RECT 2947.460 1184.490 2948.640 1185.670 ;
        RECT 2949.060 1184.490 2950.240 1185.670 ;
        RECT 2947.460 1006.090 2948.640 1007.270 ;
        RECT 2949.060 1006.090 2950.240 1007.270 ;
        RECT 2947.460 1004.490 2948.640 1005.670 ;
        RECT 2949.060 1004.490 2950.240 1005.670 ;
        RECT 2947.460 826.090 2948.640 827.270 ;
        RECT 2949.060 826.090 2950.240 827.270 ;
        RECT 2947.460 824.490 2948.640 825.670 ;
        RECT 2949.060 824.490 2950.240 825.670 ;
        RECT 2947.460 646.090 2948.640 647.270 ;
        RECT 2949.060 646.090 2950.240 647.270 ;
        RECT 2947.460 644.490 2948.640 645.670 ;
        RECT 2949.060 644.490 2950.240 645.670 ;
        RECT 2947.460 466.090 2948.640 467.270 ;
        RECT 2949.060 466.090 2950.240 467.270 ;
        RECT 2947.460 464.490 2948.640 465.670 ;
        RECT 2949.060 464.490 2950.240 465.670 ;
        RECT 2947.460 286.090 2948.640 287.270 ;
        RECT 2949.060 286.090 2950.240 287.270 ;
        RECT 2947.460 284.490 2948.640 285.670 ;
        RECT 2949.060 284.490 2950.240 285.670 ;
        RECT 2947.460 106.090 2948.640 107.270 ;
        RECT 2949.060 106.090 2950.240 107.270 ;
        RECT 2947.460 104.490 2948.640 105.670 ;
        RECT 2949.060 104.490 2950.240 105.670 ;
        RECT 2947.460 -23.660 2948.640 -22.480 ;
        RECT 2949.060 -23.660 2950.240 -22.480 ;
        RECT 2947.460 -25.260 2948.640 -24.080 ;
        RECT 2949.060 -25.260 2950.240 -24.080 ;
      LAYER met5 ;
        RECT -30.780 3542.000 2950.400 3545.100 ;
        RECT -45.180 3344.330 2964.800 3347.430 ;
        RECT -45.180 3164.330 2964.800 3167.430 ;
        RECT -45.180 2984.330 2964.800 2987.430 ;
        RECT -45.180 2804.330 2964.800 2807.430 ;
        RECT -45.180 2624.330 2964.800 2627.430 ;
        RECT -45.180 2444.330 2964.800 2447.430 ;
        RECT -45.180 2264.330 2964.800 2267.430 ;
        RECT -45.180 2084.330 2964.800 2087.430 ;
        RECT -45.180 1904.330 2964.800 1907.430 ;
        RECT -45.180 1724.330 2964.800 1727.430 ;
        RECT -45.180 1544.330 2964.800 1547.430 ;
        RECT -45.180 1364.330 2964.800 1367.430 ;
        RECT -45.180 1184.330 2964.800 1187.430 ;
        RECT -45.180 1004.330 2964.800 1007.430 ;
        RECT -45.180 824.330 2964.800 827.430 ;
        RECT -45.180 644.330 2964.800 647.430 ;
        RECT -45.180 464.330 2964.800 467.430 ;
        RECT -45.180 284.330 2964.800 287.430 ;
        RECT -45.180 104.330 2964.800 107.430 ;
        RECT -30.780 -25.420 2950.400 -22.320 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -40.380 -35.020 -37.280 3554.700 ;
        RECT 143.970 -39.820 147.070 3559.500 ;
        RECT 323.970 -39.820 327.070 3559.500 ;
        RECT 503.970 760.000 507.070 3559.500 ;
        RECT 503.970 -39.820 507.070 490.000 ;
        RECT 683.970 -39.820 687.070 3559.500 ;
        RECT 863.970 -39.820 867.070 3559.500 ;
        RECT 1043.970 -39.820 1047.070 3559.500 ;
        RECT 1223.970 -39.820 1227.070 3559.500 ;
        RECT 1403.970 -39.820 1407.070 3559.500 ;
        RECT 1583.970 -39.820 1587.070 3559.500 ;
        RECT 1763.970 -39.820 1767.070 3559.500 ;
        RECT 1943.970 -39.820 1947.070 3559.500 ;
        RECT 2123.970 -39.820 2127.070 3559.500 ;
        RECT 2303.970 -39.820 2307.070 3559.500 ;
        RECT 2483.970 -39.820 2487.070 3559.500 ;
        RECT 2663.970 -39.820 2667.070 3559.500 ;
        RECT 2843.970 -39.820 2847.070 3559.500 ;
        RECT 2956.900 -35.020 2960.000 3554.700 ;
      LAYER via4 ;
        RECT -40.220 3553.360 -39.040 3554.540 ;
        RECT -38.620 3553.360 -37.440 3554.540 ;
        RECT -40.220 3551.760 -39.040 3552.940 ;
        RECT -38.620 3551.760 -37.440 3552.940 ;
        RECT -40.220 3391.090 -39.040 3392.270 ;
        RECT -38.620 3391.090 -37.440 3392.270 ;
        RECT -40.220 3389.490 -39.040 3390.670 ;
        RECT -38.620 3389.490 -37.440 3390.670 ;
        RECT -40.220 3211.090 -39.040 3212.270 ;
        RECT -38.620 3211.090 -37.440 3212.270 ;
        RECT -40.220 3209.490 -39.040 3210.670 ;
        RECT -38.620 3209.490 -37.440 3210.670 ;
        RECT -40.220 3031.090 -39.040 3032.270 ;
        RECT -38.620 3031.090 -37.440 3032.270 ;
        RECT -40.220 3029.490 -39.040 3030.670 ;
        RECT -38.620 3029.490 -37.440 3030.670 ;
        RECT -40.220 2851.090 -39.040 2852.270 ;
        RECT -38.620 2851.090 -37.440 2852.270 ;
        RECT -40.220 2849.490 -39.040 2850.670 ;
        RECT -38.620 2849.490 -37.440 2850.670 ;
        RECT -40.220 2671.090 -39.040 2672.270 ;
        RECT -38.620 2671.090 -37.440 2672.270 ;
        RECT -40.220 2669.490 -39.040 2670.670 ;
        RECT -38.620 2669.490 -37.440 2670.670 ;
        RECT -40.220 2491.090 -39.040 2492.270 ;
        RECT -38.620 2491.090 -37.440 2492.270 ;
        RECT -40.220 2489.490 -39.040 2490.670 ;
        RECT -38.620 2489.490 -37.440 2490.670 ;
        RECT -40.220 2311.090 -39.040 2312.270 ;
        RECT -38.620 2311.090 -37.440 2312.270 ;
        RECT -40.220 2309.490 -39.040 2310.670 ;
        RECT -38.620 2309.490 -37.440 2310.670 ;
        RECT -40.220 2131.090 -39.040 2132.270 ;
        RECT -38.620 2131.090 -37.440 2132.270 ;
        RECT -40.220 2129.490 -39.040 2130.670 ;
        RECT -38.620 2129.490 -37.440 2130.670 ;
        RECT -40.220 1951.090 -39.040 1952.270 ;
        RECT -38.620 1951.090 -37.440 1952.270 ;
        RECT -40.220 1949.490 -39.040 1950.670 ;
        RECT -38.620 1949.490 -37.440 1950.670 ;
        RECT -40.220 1771.090 -39.040 1772.270 ;
        RECT -38.620 1771.090 -37.440 1772.270 ;
        RECT -40.220 1769.490 -39.040 1770.670 ;
        RECT -38.620 1769.490 -37.440 1770.670 ;
        RECT -40.220 1591.090 -39.040 1592.270 ;
        RECT -38.620 1591.090 -37.440 1592.270 ;
        RECT -40.220 1589.490 -39.040 1590.670 ;
        RECT -38.620 1589.490 -37.440 1590.670 ;
        RECT -40.220 1411.090 -39.040 1412.270 ;
        RECT -38.620 1411.090 -37.440 1412.270 ;
        RECT -40.220 1409.490 -39.040 1410.670 ;
        RECT -38.620 1409.490 -37.440 1410.670 ;
        RECT -40.220 1231.090 -39.040 1232.270 ;
        RECT -38.620 1231.090 -37.440 1232.270 ;
        RECT -40.220 1229.490 -39.040 1230.670 ;
        RECT -38.620 1229.490 -37.440 1230.670 ;
        RECT -40.220 1051.090 -39.040 1052.270 ;
        RECT -38.620 1051.090 -37.440 1052.270 ;
        RECT -40.220 1049.490 -39.040 1050.670 ;
        RECT -38.620 1049.490 -37.440 1050.670 ;
        RECT -40.220 871.090 -39.040 872.270 ;
        RECT -38.620 871.090 -37.440 872.270 ;
        RECT -40.220 869.490 -39.040 870.670 ;
        RECT -38.620 869.490 -37.440 870.670 ;
        RECT -40.220 691.090 -39.040 692.270 ;
        RECT -38.620 691.090 -37.440 692.270 ;
        RECT -40.220 689.490 -39.040 690.670 ;
        RECT -38.620 689.490 -37.440 690.670 ;
        RECT -40.220 511.090 -39.040 512.270 ;
        RECT -38.620 511.090 -37.440 512.270 ;
        RECT -40.220 509.490 -39.040 510.670 ;
        RECT -38.620 509.490 -37.440 510.670 ;
        RECT -40.220 331.090 -39.040 332.270 ;
        RECT -38.620 331.090 -37.440 332.270 ;
        RECT -40.220 329.490 -39.040 330.670 ;
        RECT -38.620 329.490 -37.440 330.670 ;
        RECT -40.220 151.090 -39.040 152.270 ;
        RECT -38.620 151.090 -37.440 152.270 ;
        RECT -40.220 149.490 -39.040 150.670 ;
        RECT -38.620 149.490 -37.440 150.670 ;
        RECT -40.220 -33.260 -39.040 -32.080 ;
        RECT -38.620 -33.260 -37.440 -32.080 ;
        RECT -40.220 -34.860 -39.040 -33.680 ;
        RECT -38.620 -34.860 -37.440 -33.680 ;
        RECT 144.130 3553.360 145.310 3554.540 ;
        RECT 145.730 3553.360 146.910 3554.540 ;
        RECT 144.130 3551.760 145.310 3552.940 ;
        RECT 145.730 3551.760 146.910 3552.940 ;
        RECT 144.130 3391.090 145.310 3392.270 ;
        RECT 145.730 3391.090 146.910 3392.270 ;
        RECT 144.130 3389.490 145.310 3390.670 ;
        RECT 145.730 3389.490 146.910 3390.670 ;
        RECT 144.130 3211.090 145.310 3212.270 ;
        RECT 145.730 3211.090 146.910 3212.270 ;
        RECT 144.130 3209.490 145.310 3210.670 ;
        RECT 145.730 3209.490 146.910 3210.670 ;
        RECT 144.130 3031.090 145.310 3032.270 ;
        RECT 145.730 3031.090 146.910 3032.270 ;
        RECT 144.130 3029.490 145.310 3030.670 ;
        RECT 145.730 3029.490 146.910 3030.670 ;
        RECT 144.130 2851.090 145.310 2852.270 ;
        RECT 145.730 2851.090 146.910 2852.270 ;
        RECT 144.130 2849.490 145.310 2850.670 ;
        RECT 145.730 2849.490 146.910 2850.670 ;
        RECT 144.130 2671.090 145.310 2672.270 ;
        RECT 145.730 2671.090 146.910 2672.270 ;
        RECT 144.130 2669.490 145.310 2670.670 ;
        RECT 145.730 2669.490 146.910 2670.670 ;
        RECT 144.130 2491.090 145.310 2492.270 ;
        RECT 145.730 2491.090 146.910 2492.270 ;
        RECT 144.130 2489.490 145.310 2490.670 ;
        RECT 145.730 2489.490 146.910 2490.670 ;
        RECT 144.130 2311.090 145.310 2312.270 ;
        RECT 145.730 2311.090 146.910 2312.270 ;
        RECT 144.130 2309.490 145.310 2310.670 ;
        RECT 145.730 2309.490 146.910 2310.670 ;
        RECT 144.130 2131.090 145.310 2132.270 ;
        RECT 145.730 2131.090 146.910 2132.270 ;
        RECT 144.130 2129.490 145.310 2130.670 ;
        RECT 145.730 2129.490 146.910 2130.670 ;
        RECT 144.130 1951.090 145.310 1952.270 ;
        RECT 145.730 1951.090 146.910 1952.270 ;
        RECT 144.130 1949.490 145.310 1950.670 ;
        RECT 145.730 1949.490 146.910 1950.670 ;
        RECT 144.130 1771.090 145.310 1772.270 ;
        RECT 145.730 1771.090 146.910 1772.270 ;
        RECT 144.130 1769.490 145.310 1770.670 ;
        RECT 145.730 1769.490 146.910 1770.670 ;
        RECT 144.130 1591.090 145.310 1592.270 ;
        RECT 145.730 1591.090 146.910 1592.270 ;
        RECT 144.130 1589.490 145.310 1590.670 ;
        RECT 145.730 1589.490 146.910 1590.670 ;
        RECT 144.130 1411.090 145.310 1412.270 ;
        RECT 145.730 1411.090 146.910 1412.270 ;
        RECT 144.130 1409.490 145.310 1410.670 ;
        RECT 145.730 1409.490 146.910 1410.670 ;
        RECT 144.130 1231.090 145.310 1232.270 ;
        RECT 145.730 1231.090 146.910 1232.270 ;
        RECT 144.130 1229.490 145.310 1230.670 ;
        RECT 145.730 1229.490 146.910 1230.670 ;
        RECT 144.130 1051.090 145.310 1052.270 ;
        RECT 145.730 1051.090 146.910 1052.270 ;
        RECT 144.130 1049.490 145.310 1050.670 ;
        RECT 145.730 1049.490 146.910 1050.670 ;
        RECT 144.130 871.090 145.310 872.270 ;
        RECT 145.730 871.090 146.910 872.270 ;
        RECT 144.130 869.490 145.310 870.670 ;
        RECT 145.730 869.490 146.910 870.670 ;
        RECT 144.130 691.090 145.310 692.270 ;
        RECT 145.730 691.090 146.910 692.270 ;
        RECT 144.130 689.490 145.310 690.670 ;
        RECT 145.730 689.490 146.910 690.670 ;
        RECT 144.130 511.090 145.310 512.270 ;
        RECT 145.730 511.090 146.910 512.270 ;
        RECT 144.130 509.490 145.310 510.670 ;
        RECT 145.730 509.490 146.910 510.670 ;
        RECT 144.130 331.090 145.310 332.270 ;
        RECT 145.730 331.090 146.910 332.270 ;
        RECT 144.130 329.490 145.310 330.670 ;
        RECT 145.730 329.490 146.910 330.670 ;
        RECT 144.130 151.090 145.310 152.270 ;
        RECT 145.730 151.090 146.910 152.270 ;
        RECT 144.130 149.490 145.310 150.670 ;
        RECT 145.730 149.490 146.910 150.670 ;
        RECT 144.130 -33.260 145.310 -32.080 ;
        RECT 145.730 -33.260 146.910 -32.080 ;
        RECT 144.130 -34.860 145.310 -33.680 ;
        RECT 145.730 -34.860 146.910 -33.680 ;
        RECT 324.130 3553.360 325.310 3554.540 ;
        RECT 325.730 3553.360 326.910 3554.540 ;
        RECT 324.130 3551.760 325.310 3552.940 ;
        RECT 325.730 3551.760 326.910 3552.940 ;
        RECT 324.130 3391.090 325.310 3392.270 ;
        RECT 325.730 3391.090 326.910 3392.270 ;
        RECT 324.130 3389.490 325.310 3390.670 ;
        RECT 325.730 3389.490 326.910 3390.670 ;
        RECT 324.130 3211.090 325.310 3212.270 ;
        RECT 325.730 3211.090 326.910 3212.270 ;
        RECT 324.130 3209.490 325.310 3210.670 ;
        RECT 325.730 3209.490 326.910 3210.670 ;
        RECT 324.130 3031.090 325.310 3032.270 ;
        RECT 325.730 3031.090 326.910 3032.270 ;
        RECT 324.130 3029.490 325.310 3030.670 ;
        RECT 325.730 3029.490 326.910 3030.670 ;
        RECT 324.130 2851.090 325.310 2852.270 ;
        RECT 325.730 2851.090 326.910 2852.270 ;
        RECT 324.130 2849.490 325.310 2850.670 ;
        RECT 325.730 2849.490 326.910 2850.670 ;
        RECT 324.130 2671.090 325.310 2672.270 ;
        RECT 325.730 2671.090 326.910 2672.270 ;
        RECT 324.130 2669.490 325.310 2670.670 ;
        RECT 325.730 2669.490 326.910 2670.670 ;
        RECT 324.130 2491.090 325.310 2492.270 ;
        RECT 325.730 2491.090 326.910 2492.270 ;
        RECT 324.130 2489.490 325.310 2490.670 ;
        RECT 325.730 2489.490 326.910 2490.670 ;
        RECT 324.130 2311.090 325.310 2312.270 ;
        RECT 325.730 2311.090 326.910 2312.270 ;
        RECT 324.130 2309.490 325.310 2310.670 ;
        RECT 325.730 2309.490 326.910 2310.670 ;
        RECT 324.130 2131.090 325.310 2132.270 ;
        RECT 325.730 2131.090 326.910 2132.270 ;
        RECT 324.130 2129.490 325.310 2130.670 ;
        RECT 325.730 2129.490 326.910 2130.670 ;
        RECT 324.130 1951.090 325.310 1952.270 ;
        RECT 325.730 1951.090 326.910 1952.270 ;
        RECT 324.130 1949.490 325.310 1950.670 ;
        RECT 325.730 1949.490 326.910 1950.670 ;
        RECT 324.130 1771.090 325.310 1772.270 ;
        RECT 325.730 1771.090 326.910 1772.270 ;
        RECT 324.130 1769.490 325.310 1770.670 ;
        RECT 325.730 1769.490 326.910 1770.670 ;
        RECT 324.130 1591.090 325.310 1592.270 ;
        RECT 325.730 1591.090 326.910 1592.270 ;
        RECT 324.130 1589.490 325.310 1590.670 ;
        RECT 325.730 1589.490 326.910 1590.670 ;
        RECT 324.130 1411.090 325.310 1412.270 ;
        RECT 325.730 1411.090 326.910 1412.270 ;
        RECT 324.130 1409.490 325.310 1410.670 ;
        RECT 325.730 1409.490 326.910 1410.670 ;
        RECT 324.130 1231.090 325.310 1232.270 ;
        RECT 325.730 1231.090 326.910 1232.270 ;
        RECT 324.130 1229.490 325.310 1230.670 ;
        RECT 325.730 1229.490 326.910 1230.670 ;
        RECT 324.130 1051.090 325.310 1052.270 ;
        RECT 325.730 1051.090 326.910 1052.270 ;
        RECT 324.130 1049.490 325.310 1050.670 ;
        RECT 325.730 1049.490 326.910 1050.670 ;
        RECT 324.130 871.090 325.310 872.270 ;
        RECT 325.730 871.090 326.910 872.270 ;
        RECT 324.130 869.490 325.310 870.670 ;
        RECT 325.730 869.490 326.910 870.670 ;
        RECT 504.130 3553.360 505.310 3554.540 ;
        RECT 505.730 3553.360 506.910 3554.540 ;
        RECT 504.130 3551.760 505.310 3552.940 ;
        RECT 505.730 3551.760 506.910 3552.940 ;
        RECT 504.130 3391.090 505.310 3392.270 ;
        RECT 505.730 3391.090 506.910 3392.270 ;
        RECT 504.130 3389.490 505.310 3390.670 ;
        RECT 505.730 3389.490 506.910 3390.670 ;
        RECT 504.130 3211.090 505.310 3212.270 ;
        RECT 505.730 3211.090 506.910 3212.270 ;
        RECT 504.130 3209.490 505.310 3210.670 ;
        RECT 505.730 3209.490 506.910 3210.670 ;
        RECT 504.130 3031.090 505.310 3032.270 ;
        RECT 505.730 3031.090 506.910 3032.270 ;
        RECT 504.130 3029.490 505.310 3030.670 ;
        RECT 505.730 3029.490 506.910 3030.670 ;
        RECT 504.130 2851.090 505.310 2852.270 ;
        RECT 505.730 2851.090 506.910 2852.270 ;
        RECT 504.130 2849.490 505.310 2850.670 ;
        RECT 505.730 2849.490 506.910 2850.670 ;
        RECT 504.130 2671.090 505.310 2672.270 ;
        RECT 505.730 2671.090 506.910 2672.270 ;
        RECT 504.130 2669.490 505.310 2670.670 ;
        RECT 505.730 2669.490 506.910 2670.670 ;
        RECT 504.130 2491.090 505.310 2492.270 ;
        RECT 505.730 2491.090 506.910 2492.270 ;
        RECT 504.130 2489.490 505.310 2490.670 ;
        RECT 505.730 2489.490 506.910 2490.670 ;
        RECT 504.130 2311.090 505.310 2312.270 ;
        RECT 505.730 2311.090 506.910 2312.270 ;
        RECT 504.130 2309.490 505.310 2310.670 ;
        RECT 505.730 2309.490 506.910 2310.670 ;
        RECT 504.130 2131.090 505.310 2132.270 ;
        RECT 505.730 2131.090 506.910 2132.270 ;
        RECT 504.130 2129.490 505.310 2130.670 ;
        RECT 505.730 2129.490 506.910 2130.670 ;
        RECT 504.130 1951.090 505.310 1952.270 ;
        RECT 505.730 1951.090 506.910 1952.270 ;
        RECT 504.130 1949.490 505.310 1950.670 ;
        RECT 505.730 1949.490 506.910 1950.670 ;
        RECT 504.130 1771.090 505.310 1772.270 ;
        RECT 505.730 1771.090 506.910 1772.270 ;
        RECT 504.130 1769.490 505.310 1770.670 ;
        RECT 505.730 1769.490 506.910 1770.670 ;
        RECT 504.130 1591.090 505.310 1592.270 ;
        RECT 505.730 1591.090 506.910 1592.270 ;
        RECT 504.130 1589.490 505.310 1590.670 ;
        RECT 505.730 1589.490 506.910 1590.670 ;
        RECT 504.130 1411.090 505.310 1412.270 ;
        RECT 505.730 1411.090 506.910 1412.270 ;
        RECT 504.130 1409.490 505.310 1410.670 ;
        RECT 505.730 1409.490 506.910 1410.670 ;
        RECT 504.130 1231.090 505.310 1232.270 ;
        RECT 505.730 1231.090 506.910 1232.270 ;
        RECT 504.130 1229.490 505.310 1230.670 ;
        RECT 505.730 1229.490 506.910 1230.670 ;
        RECT 504.130 1051.090 505.310 1052.270 ;
        RECT 505.730 1051.090 506.910 1052.270 ;
        RECT 504.130 1049.490 505.310 1050.670 ;
        RECT 505.730 1049.490 506.910 1050.670 ;
        RECT 504.130 871.090 505.310 872.270 ;
        RECT 505.730 871.090 506.910 872.270 ;
        RECT 504.130 869.490 505.310 870.670 ;
        RECT 505.730 869.490 506.910 870.670 ;
        RECT 684.130 3553.360 685.310 3554.540 ;
        RECT 685.730 3553.360 686.910 3554.540 ;
        RECT 684.130 3551.760 685.310 3552.940 ;
        RECT 685.730 3551.760 686.910 3552.940 ;
        RECT 684.130 3391.090 685.310 3392.270 ;
        RECT 685.730 3391.090 686.910 3392.270 ;
        RECT 684.130 3389.490 685.310 3390.670 ;
        RECT 685.730 3389.490 686.910 3390.670 ;
        RECT 684.130 3211.090 685.310 3212.270 ;
        RECT 685.730 3211.090 686.910 3212.270 ;
        RECT 684.130 3209.490 685.310 3210.670 ;
        RECT 685.730 3209.490 686.910 3210.670 ;
        RECT 684.130 3031.090 685.310 3032.270 ;
        RECT 685.730 3031.090 686.910 3032.270 ;
        RECT 684.130 3029.490 685.310 3030.670 ;
        RECT 685.730 3029.490 686.910 3030.670 ;
        RECT 684.130 2851.090 685.310 2852.270 ;
        RECT 685.730 2851.090 686.910 2852.270 ;
        RECT 684.130 2849.490 685.310 2850.670 ;
        RECT 685.730 2849.490 686.910 2850.670 ;
        RECT 684.130 2671.090 685.310 2672.270 ;
        RECT 685.730 2671.090 686.910 2672.270 ;
        RECT 684.130 2669.490 685.310 2670.670 ;
        RECT 685.730 2669.490 686.910 2670.670 ;
        RECT 684.130 2491.090 685.310 2492.270 ;
        RECT 685.730 2491.090 686.910 2492.270 ;
        RECT 684.130 2489.490 685.310 2490.670 ;
        RECT 685.730 2489.490 686.910 2490.670 ;
        RECT 684.130 2311.090 685.310 2312.270 ;
        RECT 685.730 2311.090 686.910 2312.270 ;
        RECT 684.130 2309.490 685.310 2310.670 ;
        RECT 685.730 2309.490 686.910 2310.670 ;
        RECT 684.130 2131.090 685.310 2132.270 ;
        RECT 685.730 2131.090 686.910 2132.270 ;
        RECT 684.130 2129.490 685.310 2130.670 ;
        RECT 685.730 2129.490 686.910 2130.670 ;
        RECT 684.130 1951.090 685.310 1952.270 ;
        RECT 685.730 1951.090 686.910 1952.270 ;
        RECT 684.130 1949.490 685.310 1950.670 ;
        RECT 685.730 1949.490 686.910 1950.670 ;
        RECT 684.130 1771.090 685.310 1772.270 ;
        RECT 685.730 1771.090 686.910 1772.270 ;
        RECT 684.130 1769.490 685.310 1770.670 ;
        RECT 685.730 1769.490 686.910 1770.670 ;
        RECT 684.130 1591.090 685.310 1592.270 ;
        RECT 685.730 1591.090 686.910 1592.270 ;
        RECT 684.130 1589.490 685.310 1590.670 ;
        RECT 685.730 1589.490 686.910 1590.670 ;
        RECT 684.130 1411.090 685.310 1412.270 ;
        RECT 685.730 1411.090 686.910 1412.270 ;
        RECT 684.130 1409.490 685.310 1410.670 ;
        RECT 685.730 1409.490 686.910 1410.670 ;
        RECT 684.130 1231.090 685.310 1232.270 ;
        RECT 685.730 1231.090 686.910 1232.270 ;
        RECT 684.130 1229.490 685.310 1230.670 ;
        RECT 685.730 1229.490 686.910 1230.670 ;
        RECT 684.130 1051.090 685.310 1052.270 ;
        RECT 685.730 1051.090 686.910 1052.270 ;
        RECT 684.130 1049.490 685.310 1050.670 ;
        RECT 685.730 1049.490 686.910 1050.670 ;
        RECT 684.130 871.090 685.310 872.270 ;
        RECT 685.730 871.090 686.910 872.270 ;
        RECT 684.130 869.490 685.310 870.670 ;
        RECT 685.730 869.490 686.910 870.670 ;
        RECT 324.130 691.090 325.310 692.270 ;
        RECT 325.730 691.090 326.910 692.270 ;
        RECT 324.130 689.490 325.310 690.670 ;
        RECT 325.730 689.490 326.910 690.670 ;
        RECT 324.130 511.090 325.310 512.270 ;
        RECT 325.730 511.090 326.910 512.270 ;
        RECT 324.130 509.490 325.310 510.670 ;
        RECT 325.730 509.490 326.910 510.670 ;
        RECT 684.130 691.090 685.310 692.270 ;
        RECT 685.730 691.090 686.910 692.270 ;
        RECT 684.130 689.490 685.310 690.670 ;
        RECT 685.730 689.490 686.910 690.670 ;
        RECT 684.130 511.090 685.310 512.270 ;
        RECT 685.730 511.090 686.910 512.270 ;
        RECT 684.130 509.490 685.310 510.670 ;
        RECT 685.730 509.490 686.910 510.670 ;
        RECT 324.130 331.090 325.310 332.270 ;
        RECT 325.730 331.090 326.910 332.270 ;
        RECT 324.130 329.490 325.310 330.670 ;
        RECT 325.730 329.490 326.910 330.670 ;
        RECT 324.130 151.090 325.310 152.270 ;
        RECT 325.730 151.090 326.910 152.270 ;
        RECT 324.130 149.490 325.310 150.670 ;
        RECT 325.730 149.490 326.910 150.670 ;
        RECT 324.130 -33.260 325.310 -32.080 ;
        RECT 325.730 -33.260 326.910 -32.080 ;
        RECT 324.130 -34.860 325.310 -33.680 ;
        RECT 325.730 -34.860 326.910 -33.680 ;
        RECT 504.130 331.090 505.310 332.270 ;
        RECT 505.730 331.090 506.910 332.270 ;
        RECT 504.130 329.490 505.310 330.670 ;
        RECT 505.730 329.490 506.910 330.670 ;
        RECT 504.130 151.090 505.310 152.270 ;
        RECT 505.730 151.090 506.910 152.270 ;
        RECT 504.130 149.490 505.310 150.670 ;
        RECT 505.730 149.490 506.910 150.670 ;
        RECT 504.130 -33.260 505.310 -32.080 ;
        RECT 505.730 -33.260 506.910 -32.080 ;
        RECT 504.130 -34.860 505.310 -33.680 ;
        RECT 505.730 -34.860 506.910 -33.680 ;
        RECT 684.130 331.090 685.310 332.270 ;
        RECT 685.730 331.090 686.910 332.270 ;
        RECT 684.130 329.490 685.310 330.670 ;
        RECT 685.730 329.490 686.910 330.670 ;
        RECT 684.130 151.090 685.310 152.270 ;
        RECT 685.730 151.090 686.910 152.270 ;
        RECT 684.130 149.490 685.310 150.670 ;
        RECT 685.730 149.490 686.910 150.670 ;
        RECT 684.130 -33.260 685.310 -32.080 ;
        RECT 685.730 -33.260 686.910 -32.080 ;
        RECT 684.130 -34.860 685.310 -33.680 ;
        RECT 685.730 -34.860 686.910 -33.680 ;
        RECT 864.130 3553.360 865.310 3554.540 ;
        RECT 865.730 3553.360 866.910 3554.540 ;
        RECT 864.130 3551.760 865.310 3552.940 ;
        RECT 865.730 3551.760 866.910 3552.940 ;
        RECT 864.130 3391.090 865.310 3392.270 ;
        RECT 865.730 3391.090 866.910 3392.270 ;
        RECT 864.130 3389.490 865.310 3390.670 ;
        RECT 865.730 3389.490 866.910 3390.670 ;
        RECT 864.130 3211.090 865.310 3212.270 ;
        RECT 865.730 3211.090 866.910 3212.270 ;
        RECT 864.130 3209.490 865.310 3210.670 ;
        RECT 865.730 3209.490 866.910 3210.670 ;
        RECT 864.130 3031.090 865.310 3032.270 ;
        RECT 865.730 3031.090 866.910 3032.270 ;
        RECT 864.130 3029.490 865.310 3030.670 ;
        RECT 865.730 3029.490 866.910 3030.670 ;
        RECT 864.130 2851.090 865.310 2852.270 ;
        RECT 865.730 2851.090 866.910 2852.270 ;
        RECT 864.130 2849.490 865.310 2850.670 ;
        RECT 865.730 2849.490 866.910 2850.670 ;
        RECT 864.130 2671.090 865.310 2672.270 ;
        RECT 865.730 2671.090 866.910 2672.270 ;
        RECT 864.130 2669.490 865.310 2670.670 ;
        RECT 865.730 2669.490 866.910 2670.670 ;
        RECT 864.130 2491.090 865.310 2492.270 ;
        RECT 865.730 2491.090 866.910 2492.270 ;
        RECT 864.130 2489.490 865.310 2490.670 ;
        RECT 865.730 2489.490 866.910 2490.670 ;
        RECT 864.130 2311.090 865.310 2312.270 ;
        RECT 865.730 2311.090 866.910 2312.270 ;
        RECT 864.130 2309.490 865.310 2310.670 ;
        RECT 865.730 2309.490 866.910 2310.670 ;
        RECT 864.130 2131.090 865.310 2132.270 ;
        RECT 865.730 2131.090 866.910 2132.270 ;
        RECT 864.130 2129.490 865.310 2130.670 ;
        RECT 865.730 2129.490 866.910 2130.670 ;
        RECT 864.130 1951.090 865.310 1952.270 ;
        RECT 865.730 1951.090 866.910 1952.270 ;
        RECT 864.130 1949.490 865.310 1950.670 ;
        RECT 865.730 1949.490 866.910 1950.670 ;
        RECT 864.130 1771.090 865.310 1772.270 ;
        RECT 865.730 1771.090 866.910 1772.270 ;
        RECT 864.130 1769.490 865.310 1770.670 ;
        RECT 865.730 1769.490 866.910 1770.670 ;
        RECT 864.130 1591.090 865.310 1592.270 ;
        RECT 865.730 1591.090 866.910 1592.270 ;
        RECT 864.130 1589.490 865.310 1590.670 ;
        RECT 865.730 1589.490 866.910 1590.670 ;
        RECT 864.130 1411.090 865.310 1412.270 ;
        RECT 865.730 1411.090 866.910 1412.270 ;
        RECT 864.130 1409.490 865.310 1410.670 ;
        RECT 865.730 1409.490 866.910 1410.670 ;
        RECT 864.130 1231.090 865.310 1232.270 ;
        RECT 865.730 1231.090 866.910 1232.270 ;
        RECT 864.130 1229.490 865.310 1230.670 ;
        RECT 865.730 1229.490 866.910 1230.670 ;
        RECT 864.130 1051.090 865.310 1052.270 ;
        RECT 865.730 1051.090 866.910 1052.270 ;
        RECT 864.130 1049.490 865.310 1050.670 ;
        RECT 865.730 1049.490 866.910 1050.670 ;
        RECT 864.130 871.090 865.310 872.270 ;
        RECT 865.730 871.090 866.910 872.270 ;
        RECT 864.130 869.490 865.310 870.670 ;
        RECT 865.730 869.490 866.910 870.670 ;
        RECT 864.130 691.090 865.310 692.270 ;
        RECT 865.730 691.090 866.910 692.270 ;
        RECT 864.130 689.490 865.310 690.670 ;
        RECT 865.730 689.490 866.910 690.670 ;
        RECT 864.130 511.090 865.310 512.270 ;
        RECT 865.730 511.090 866.910 512.270 ;
        RECT 864.130 509.490 865.310 510.670 ;
        RECT 865.730 509.490 866.910 510.670 ;
        RECT 864.130 331.090 865.310 332.270 ;
        RECT 865.730 331.090 866.910 332.270 ;
        RECT 864.130 329.490 865.310 330.670 ;
        RECT 865.730 329.490 866.910 330.670 ;
        RECT 864.130 151.090 865.310 152.270 ;
        RECT 865.730 151.090 866.910 152.270 ;
        RECT 864.130 149.490 865.310 150.670 ;
        RECT 865.730 149.490 866.910 150.670 ;
        RECT 864.130 -33.260 865.310 -32.080 ;
        RECT 865.730 -33.260 866.910 -32.080 ;
        RECT 864.130 -34.860 865.310 -33.680 ;
        RECT 865.730 -34.860 866.910 -33.680 ;
        RECT 1044.130 3553.360 1045.310 3554.540 ;
        RECT 1045.730 3553.360 1046.910 3554.540 ;
        RECT 1044.130 3551.760 1045.310 3552.940 ;
        RECT 1045.730 3551.760 1046.910 3552.940 ;
        RECT 1044.130 3391.090 1045.310 3392.270 ;
        RECT 1045.730 3391.090 1046.910 3392.270 ;
        RECT 1044.130 3389.490 1045.310 3390.670 ;
        RECT 1045.730 3389.490 1046.910 3390.670 ;
        RECT 1044.130 3211.090 1045.310 3212.270 ;
        RECT 1045.730 3211.090 1046.910 3212.270 ;
        RECT 1044.130 3209.490 1045.310 3210.670 ;
        RECT 1045.730 3209.490 1046.910 3210.670 ;
        RECT 1044.130 3031.090 1045.310 3032.270 ;
        RECT 1045.730 3031.090 1046.910 3032.270 ;
        RECT 1044.130 3029.490 1045.310 3030.670 ;
        RECT 1045.730 3029.490 1046.910 3030.670 ;
        RECT 1044.130 2851.090 1045.310 2852.270 ;
        RECT 1045.730 2851.090 1046.910 2852.270 ;
        RECT 1044.130 2849.490 1045.310 2850.670 ;
        RECT 1045.730 2849.490 1046.910 2850.670 ;
        RECT 1044.130 2671.090 1045.310 2672.270 ;
        RECT 1045.730 2671.090 1046.910 2672.270 ;
        RECT 1044.130 2669.490 1045.310 2670.670 ;
        RECT 1045.730 2669.490 1046.910 2670.670 ;
        RECT 1044.130 2491.090 1045.310 2492.270 ;
        RECT 1045.730 2491.090 1046.910 2492.270 ;
        RECT 1044.130 2489.490 1045.310 2490.670 ;
        RECT 1045.730 2489.490 1046.910 2490.670 ;
        RECT 1044.130 2311.090 1045.310 2312.270 ;
        RECT 1045.730 2311.090 1046.910 2312.270 ;
        RECT 1044.130 2309.490 1045.310 2310.670 ;
        RECT 1045.730 2309.490 1046.910 2310.670 ;
        RECT 1044.130 2131.090 1045.310 2132.270 ;
        RECT 1045.730 2131.090 1046.910 2132.270 ;
        RECT 1044.130 2129.490 1045.310 2130.670 ;
        RECT 1045.730 2129.490 1046.910 2130.670 ;
        RECT 1044.130 1951.090 1045.310 1952.270 ;
        RECT 1045.730 1951.090 1046.910 1952.270 ;
        RECT 1044.130 1949.490 1045.310 1950.670 ;
        RECT 1045.730 1949.490 1046.910 1950.670 ;
        RECT 1044.130 1771.090 1045.310 1772.270 ;
        RECT 1045.730 1771.090 1046.910 1772.270 ;
        RECT 1044.130 1769.490 1045.310 1770.670 ;
        RECT 1045.730 1769.490 1046.910 1770.670 ;
        RECT 1044.130 1591.090 1045.310 1592.270 ;
        RECT 1045.730 1591.090 1046.910 1592.270 ;
        RECT 1044.130 1589.490 1045.310 1590.670 ;
        RECT 1045.730 1589.490 1046.910 1590.670 ;
        RECT 1044.130 1411.090 1045.310 1412.270 ;
        RECT 1045.730 1411.090 1046.910 1412.270 ;
        RECT 1044.130 1409.490 1045.310 1410.670 ;
        RECT 1045.730 1409.490 1046.910 1410.670 ;
        RECT 1044.130 1231.090 1045.310 1232.270 ;
        RECT 1045.730 1231.090 1046.910 1232.270 ;
        RECT 1044.130 1229.490 1045.310 1230.670 ;
        RECT 1045.730 1229.490 1046.910 1230.670 ;
        RECT 1044.130 1051.090 1045.310 1052.270 ;
        RECT 1045.730 1051.090 1046.910 1052.270 ;
        RECT 1044.130 1049.490 1045.310 1050.670 ;
        RECT 1045.730 1049.490 1046.910 1050.670 ;
        RECT 1044.130 871.090 1045.310 872.270 ;
        RECT 1045.730 871.090 1046.910 872.270 ;
        RECT 1044.130 869.490 1045.310 870.670 ;
        RECT 1045.730 869.490 1046.910 870.670 ;
        RECT 1044.130 691.090 1045.310 692.270 ;
        RECT 1045.730 691.090 1046.910 692.270 ;
        RECT 1044.130 689.490 1045.310 690.670 ;
        RECT 1045.730 689.490 1046.910 690.670 ;
        RECT 1044.130 511.090 1045.310 512.270 ;
        RECT 1045.730 511.090 1046.910 512.270 ;
        RECT 1044.130 509.490 1045.310 510.670 ;
        RECT 1045.730 509.490 1046.910 510.670 ;
        RECT 1044.130 331.090 1045.310 332.270 ;
        RECT 1045.730 331.090 1046.910 332.270 ;
        RECT 1044.130 329.490 1045.310 330.670 ;
        RECT 1045.730 329.490 1046.910 330.670 ;
        RECT 1044.130 151.090 1045.310 152.270 ;
        RECT 1045.730 151.090 1046.910 152.270 ;
        RECT 1044.130 149.490 1045.310 150.670 ;
        RECT 1045.730 149.490 1046.910 150.670 ;
        RECT 1044.130 -33.260 1045.310 -32.080 ;
        RECT 1045.730 -33.260 1046.910 -32.080 ;
        RECT 1044.130 -34.860 1045.310 -33.680 ;
        RECT 1045.730 -34.860 1046.910 -33.680 ;
        RECT 1224.130 3553.360 1225.310 3554.540 ;
        RECT 1225.730 3553.360 1226.910 3554.540 ;
        RECT 1224.130 3551.760 1225.310 3552.940 ;
        RECT 1225.730 3551.760 1226.910 3552.940 ;
        RECT 1224.130 3391.090 1225.310 3392.270 ;
        RECT 1225.730 3391.090 1226.910 3392.270 ;
        RECT 1224.130 3389.490 1225.310 3390.670 ;
        RECT 1225.730 3389.490 1226.910 3390.670 ;
        RECT 1224.130 3211.090 1225.310 3212.270 ;
        RECT 1225.730 3211.090 1226.910 3212.270 ;
        RECT 1224.130 3209.490 1225.310 3210.670 ;
        RECT 1225.730 3209.490 1226.910 3210.670 ;
        RECT 1224.130 3031.090 1225.310 3032.270 ;
        RECT 1225.730 3031.090 1226.910 3032.270 ;
        RECT 1224.130 3029.490 1225.310 3030.670 ;
        RECT 1225.730 3029.490 1226.910 3030.670 ;
        RECT 1224.130 2851.090 1225.310 2852.270 ;
        RECT 1225.730 2851.090 1226.910 2852.270 ;
        RECT 1224.130 2849.490 1225.310 2850.670 ;
        RECT 1225.730 2849.490 1226.910 2850.670 ;
        RECT 1224.130 2671.090 1225.310 2672.270 ;
        RECT 1225.730 2671.090 1226.910 2672.270 ;
        RECT 1224.130 2669.490 1225.310 2670.670 ;
        RECT 1225.730 2669.490 1226.910 2670.670 ;
        RECT 1224.130 2491.090 1225.310 2492.270 ;
        RECT 1225.730 2491.090 1226.910 2492.270 ;
        RECT 1224.130 2489.490 1225.310 2490.670 ;
        RECT 1225.730 2489.490 1226.910 2490.670 ;
        RECT 1224.130 2311.090 1225.310 2312.270 ;
        RECT 1225.730 2311.090 1226.910 2312.270 ;
        RECT 1224.130 2309.490 1225.310 2310.670 ;
        RECT 1225.730 2309.490 1226.910 2310.670 ;
        RECT 1224.130 2131.090 1225.310 2132.270 ;
        RECT 1225.730 2131.090 1226.910 2132.270 ;
        RECT 1224.130 2129.490 1225.310 2130.670 ;
        RECT 1225.730 2129.490 1226.910 2130.670 ;
        RECT 1224.130 1951.090 1225.310 1952.270 ;
        RECT 1225.730 1951.090 1226.910 1952.270 ;
        RECT 1224.130 1949.490 1225.310 1950.670 ;
        RECT 1225.730 1949.490 1226.910 1950.670 ;
        RECT 1224.130 1771.090 1225.310 1772.270 ;
        RECT 1225.730 1771.090 1226.910 1772.270 ;
        RECT 1224.130 1769.490 1225.310 1770.670 ;
        RECT 1225.730 1769.490 1226.910 1770.670 ;
        RECT 1224.130 1591.090 1225.310 1592.270 ;
        RECT 1225.730 1591.090 1226.910 1592.270 ;
        RECT 1224.130 1589.490 1225.310 1590.670 ;
        RECT 1225.730 1589.490 1226.910 1590.670 ;
        RECT 1224.130 1411.090 1225.310 1412.270 ;
        RECT 1225.730 1411.090 1226.910 1412.270 ;
        RECT 1224.130 1409.490 1225.310 1410.670 ;
        RECT 1225.730 1409.490 1226.910 1410.670 ;
        RECT 1224.130 1231.090 1225.310 1232.270 ;
        RECT 1225.730 1231.090 1226.910 1232.270 ;
        RECT 1224.130 1229.490 1225.310 1230.670 ;
        RECT 1225.730 1229.490 1226.910 1230.670 ;
        RECT 1224.130 1051.090 1225.310 1052.270 ;
        RECT 1225.730 1051.090 1226.910 1052.270 ;
        RECT 1224.130 1049.490 1225.310 1050.670 ;
        RECT 1225.730 1049.490 1226.910 1050.670 ;
        RECT 1224.130 871.090 1225.310 872.270 ;
        RECT 1225.730 871.090 1226.910 872.270 ;
        RECT 1224.130 869.490 1225.310 870.670 ;
        RECT 1225.730 869.490 1226.910 870.670 ;
        RECT 1224.130 691.090 1225.310 692.270 ;
        RECT 1225.730 691.090 1226.910 692.270 ;
        RECT 1224.130 689.490 1225.310 690.670 ;
        RECT 1225.730 689.490 1226.910 690.670 ;
        RECT 1224.130 511.090 1225.310 512.270 ;
        RECT 1225.730 511.090 1226.910 512.270 ;
        RECT 1224.130 509.490 1225.310 510.670 ;
        RECT 1225.730 509.490 1226.910 510.670 ;
        RECT 1224.130 331.090 1225.310 332.270 ;
        RECT 1225.730 331.090 1226.910 332.270 ;
        RECT 1224.130 329.490 1225.310 330.670 ;
        RECT 1225.730 329.490 1226.910 330.670 ;
        RECT 1224.130 151.090 1225.310 152.270 ;
        RECT 1225.730 151.090 1226.910 152.270 ;
        RECT 1224.130 149.490 1225.310 150.670 ;
        RECT 1225.730 149.490 1226.910 150.670 ;
        RECT 1224.130 -33.260 1225.310 -32.080 ;
        RECT 1225.730 -33.260 1226.910 -32.080 ;
        RECT 1224.130 -34.860 1225.310 -33.680 ;
        RECT 1225.730 -34.860 1226.910 -33.680 ;
        RECT 1404.130 3553.360 1405.310 3554.540 ;
        RECT 1405.730 3553.360 1406.910 3554.540 ;
        RECT 1404.130 3551.760 1405.310 3552.940 ;
        RECT 1405.730 3551.760 1406.910 3552.940 ;
        RECT 1404.130 3391.090 1405.310 3392.270 ;
        RECT 1405.730 3391.090 1406.910 3392.270 ;
        RECT 1404.130 3389.490 1405.310 3390.670 ;
        RECT 1405.730 3389.490 1406.910 3390.670 ;
        RECT 1404.130 3211.090 1405.310 3212.270 ;
        RECT 1405.730 3211.090 1406.910 3212.270 ;
        RECT 1404.130 3209.490 1405.310 3210.670 ;
        RECT 1405.730 3209.490 1406.910 3210.670 ;
        RECT 1404.130 3031.090 1405.310 3032.270 ;
        RECT 1405.730 3031.090 1406.910 3032.270 ;
        RECT 1404.130 3029.490 1405.310 3030.670 ;
        RECT 1405.730 3029.490 1406.910 3030.670 ;
        RECT 1404.130 2851.090 1405.310 2852.270 ;
        RECT 1405.730 2851.090 1406.910 2852.270 ;
        RECT 1404.130 2849.490 1405.310 2850.670 ;
        RECT 1405.730 2849.490 1406.910 2850.670 ;
        RECT 1404.130 2671.090 1405.310 2672.270 ;
        RECT 1405.730 2671.090 1406.910 2672.270 ;
        RECT 1404.130 2669.490 1405.310 2670.670 ;
        RECT 1405.730 2669.490 1406.910 2670.670 ;
        RECT 1404.130 2491.090 1405.310 2492.270 ;
        RECT 1405.730 2491.090 1406.910 2492.270 ;
        RECT 1404.130 2489.490 1405.310 2490.670 ;
        RECT 1405.730 2489.490 1406.910 2490.670 ;
        RECT 1404.130 2311.090 1405.310 2312.270 ;
        RECT 1405.730 2311.090 1406.910 2312.270 ;
        RECT 1404.130 2309.490 1405.310 2310.670 ;
        RECT 1405.730 2309.490 1406.910 2310.670 ;
        RECT 1404.130 2131.090 1405.310 2132.270 ;
        RECT 1405.730 2131.090 1406.910 2132.270 ;
        RECT 1404.130 2129.490 1405.310 2130.670 ;
        RECT 1405.730 2129.490 1406.910 2130.670 ;
        RECT 1404.130 1951.090 1405.310 1952.270 ;
        RECT 1405.730 1951.090 1406.910 1952.270 ;
        RECT 1404.130 1949.490 1405.310 1950.670 ;
        RECT 1405.730 1949.490 1406.910 1950.670 ;
        RECT 1404.130 1771.090 1405.310 1772.270 ;
        RECT 1405.730 1771.090 1406.910 1772.270 ;
        RECT 1404.130 1769.490 1405.310 1770.670 ;
        RECT 1405.730 1769.490 1406.910 1770.670 ;
        RECT 1404.130 1591.090 1405.310 1592.270 ;
        RECT 1405.730 1591.090 1406.910 1592.270 ;
        RECT 1404.130 1589.490 1405.310 1590.670 ;
        RECT 1405.730 1589.490 1406.910 1590.670 ;
        RECT 1404.130 1411.090 1405.310 1412.270 ;
        RECT 1405.730 1411.090 1406.910 1412.270 ;
        RECT 1404.130 1409.490 1405.310 1410.670 ;
        RECT 1405.730 1409.490 1406.910 1410.670 ;
        RECT 1404.130 1231.090 1405.310 1232.270 ;
        RECT 1405.730 1231.090 1406.910 1232.270 ;
        RECT 1404.130 1229.490 1405.310 1230.670 ;
        RECT 1405.730 1229.490 1406.910 1230.670 ;
        RECT 1404.130 1051.090 1405.310 1052.270 ;
        RECT 1405.730 1051.090 1406.910 1052.270 ;
        RECT 1404.130 1049.490 1405.310 1050.670 ;
        RECT 1405.730 1049.490 1406.910 1050.670 ;
        RECT 1404.130 871.090 1405.310 872.270 ;
        RECT 1405.730 871.090 1406.910 872.270 ;
        RECT 1404.130 869.490 1405.310 870.670 ;
        RECT 1405.730 869.490 1406.910 870.670 ;
        RECT 1404.130 691.090 1405.310 692.270 ;
        RECT 1405.730 691.090 1406.910 692.270 ;
        RECT 1404.130 689.490 1405.310 690.670 ;
        RECT 1405.730 689.490 1406.910 690.670 ;
        RECT 1404.130 511.090 1405.310 512.270 ;
        RECT 1405.730 511.090 1406.910 512.270 ;
        RECT 1404.130 509.490 1405.310 510.670 ;
        RECT 1405.730 509.490 1406.910 510.670 ;
        RECT 1404.130 331.090 1405.310 332.270 ;
        RECT 1405.730 331.090 1406.910 332.270 ;
        RECT 1404.130 329.490 1405.310 330.670 ;
        RECT 1405.730 329.490 1406.910 330.670 ;
        RECT 1404.130 151.090 1405.310 152.270 ;
        RECT 1405.730 151.090 1406.910 152.270 ;
        RECT 1404.130 149.490 1405.310 150.670 ;
        RECT 1405.730 149.490 1406.910 150.670 ;
        RECT 1404.130 -33.260 1405.310 -32.080 ;
        RECT 1405.730 -33.260 1406.910 -32.080 ;
        RECT 1404.130 -34.860 1405.310 -33.680 ;
        RECT 1405.730 -34.860 1406.910 -33.680 ;
        RECT 1584.130 3553.360 1585.310 3554.540 ;
        RECT 1585.730 3553.360 1586.910 3554.540 ;
        RECT 1584.130 3551.760 1585.310 3552.940 ;
        RECT 1585.730 3551.760 1586.910 3552.940 ;
        RECT 1584.130 3391.090 1585.310 3392.270 ;
        RECT 1585.730 3391.090 1586.910 3392.270 ;
        RECT 1584.130 3389.490 1585.310 3390.670 ;
        RECT 1585.730 3389.490 1586.910 3390.670 ;
        RECT 1584.130 3211.090 1585.310 3212.270 ;
        RECT 1585.730 3211.090 1586.910 3212.270 ;
        RECT 1584.130 3209.490 1585.310 3210.670 ;
        RECT 1585.730 3209.490 1586.910 3210.670 ;
        RECT 1584.130 3031.090 1585.310 3032.270 ;
        RECT 1585.730 3031.090 1586.910 3032.270 ;
        RECT 1584.130 3029.490 1585.310 3030.670 ;
        RECT 1585.730 3029.490 1586.910 3030.670 ;
        RECT 1584.130 2851.090 1585.310 2852.270 ;
        RECT 1585.730 2851.090 1586.910 2852.270 ;
        RECT 1584.130 2849.490 1585.310 2850.670 ;
        RECT 1585.730 2849.490 1586.910 2850.670 ;
        RECT 1584.130 2671.090 1585.310 2672.270 ;
        RECT 1585.730 2671.090 1586.910 2672.270 ;
        RECT 1584.130 2669.490 1585.310 2670.670 ;
        RECT 1585.730 2669.490 1586.910 2670.670 ;
        RECT 1584.130 2491.090 1585.310 2492.270 ;
        RECT 1585.730 2491.090 1586.910 2492.270 ;
        RECT 1584.130 2489.490 1585.310 2490.670 ;
        RECT 1585.730 2489.490 1586.910 2490.670 ;
        RECT 1584.130 2311.090 1585.310 2312.270 ;
        RECT 1585.730 2311.090 1586.910 2312.270 ;
        RECT 1584.130 2309.490 1585.310 2310.670 ;
        RECT 1585.730 2309.490 1586.910 2310.670 ;
        RECT 1584.130 2131.090 1585.310 2132.270 ;
        RECT 1585.730 2131.090 1586.910 2132.270 ;
        RECT 1584.130 2129.490 1585.310 2130.670 ;
        RECT 1585.730 2129.490 1586.910 2130.670 ;
        RECT 1584.130 1951.090 1585.310 1952.270 ;
        RECT 1585.730 1951.090 1586.910 1952.270 ;
        RECT 1584.130 1949.490 1585.310 1950.670 ;
        RECT 1585.730 1949.490 1586.910 1950.670 ;
        RECT 1584.130 1771.090 1585.310 1772.270 ;
        RECT 1585.730 1771.090 1586.910 1772.270 ;
        RECT 1584.130 1769.490 1585.310 1770.670 ;
        RECT 1585.730 1769.490 1586.910 1770.670 ;
        RECT 1584.130 1591.090 1585.310 1592.270 ;
        RECT 1585.730 1591.090 1586.910 1592.270 ;
        RECT 1584.130 1589.490 1585.310 1590.670 ;
        RECT 1585.730 1589.490 1586.910 1590.670 ;
        RECT 1584.130 1411.090 1585.310 1412.270 ;
        RECT 1585.730 1411.090 1586.910 1412.270 ;
        RECT 1584.130 1409.490 1585.310 1410.670 ;
        RECT 1585.730 1409.490 1586.910 1410.670 ;
        RECT 1584.130 1231.090 1585.310 1232.270 ;
        RECT 1585.730 1231.090 1586.910 1232.270 ;
        RECT 1584.130 1229.490 1585.310 1230.670 ;
        RECT 1585.730 1229.490 1586.910 1230.670 ;
        RECT 1584.130 1051.090 1585.310 1052.270 ;
        RECT 1585.730 1051.090 1586.910 1052.270 ;
        RECT 1584.130 1049.490 1585.310 1050.670 ;
        RECT 1585.730 1049.490 1586.910 1050.670 ;
        RECT 1584.130 871.090 1585.310 872.270 ;
        RECT 1585.730 871.090 1586.910 872.270 ;
        RECT 1584.130 869.490 1585.310 870.670 ;
        RECT 1585.730 869.490 1586.910 870.670 ;
        RECT 1584.130 691.090 1585.310 692.270 ;
        RECT 1585.730 691.090 1586.910 692.270 ;
        RECT 1584.130 689.490 1585.310 690.670 ;
        RECT 1585.730 689.490 1586.910 690.670 ;
        RECT 1584.130 511.090 1585.310 512.270 ;
        RECT 1585.730 511.090 1586.910 512.270 ;
        RECT 1584.130 509.490 1585.310 510.670 ;
        RECT 1585.730 509.490 1586.910 510.670 ;
        RECT 1584.130 331.090 1585.310 332.270 ;
        RECT 1585.730 331.090 1586.910 332.270 ;
        RECT 1584.130 329.490 1585.310 330.670 ;
        RECT 1585.730 329.490 1586.910 330.670 ;
        RECT 1584.130 151.090 1585.310 152.270 ;
        RECT 1585.730 151.090 1586.910 152.270 ;
        RECT 1584.130 149.490 1585.310 150.670 ;
        RECT 1585.730 149.490 1586.910 150.670 ;
        RECT 1584.130 -33.260 1585.310 -32.080 ;
        RECT 1585.730 -33.260 1586.910 -32.080 ;
        RECT 1584.130 -34.860 1585.310 -33.680 ;
        RECT 1585.730 -34.860 1586.910 -33.680 ;
        RECT 1764.130 3553.360 1765.310 3554.540 ;
        RECT 1765.730 3553.360 1766.910 3554.540 ;
        RECT 1764.130 3551.760 1765.310 3552.940 ;
        RECT 1765.730 3551.760 1766.910 3552.940 ;
        RECT 1764.130 3391.090 1765.310 3392.270 ;
        RECT 1765.730 3391.090 1766.910 3392.270 ;
        RECT 1764.130 3389.490 1765.310 3390.670 ;
        RECT 1765.730 3389.490 1766.910 3390.670 ;
        RECT 1764.130 3211.090 1765.310 3212.270 ;
        RECT 1765.730 3211.090 1766.910 3212.270 ;
        RECT 1764.130 3209.490 1765.310 3210.670 ;
        RECT 1765.730 3209.490 1766.910 3210.670 ;
        RECT 1764.130 3031.090 1765.310 3032.270 ;
        RECT 1765.730 3031.090 1766.910 3032.270 ;
        RECT 1764.130 3029.490 1765.310 3030.670 ;
        RECT 1765.730 3029.490 1766.910 3030.670 ;
        RECT 1764.130 2851.090 1765.310 2852.270 ;
        RECT 1765.730 2851.090 1766.910 2852.270 ;
        RECT 1764.130 2849.490 1765.310 2850.670 ;
        RECT 1765.730 2849.490 1766.910 2850.670 ;
        RECT 1764.130 2671.090 1765.310 2672.270 ;
        RECT 1765.730 2671.090 1766.910 2672.270 ;
        RECT 1764.130 2669.490 1765.310 2670.670 ;
        RECT 1765.730 2669.490 1766.910 2670.670 ;
        RECT 1764.130 2491.090 1765.310 2492.270 ;
        RECT 1765.730 2491.090 1766.910 2492.270 ;
        RECT 1764.130 2489.490 1765.310 2490.670 ;
        RECT 1765.730 2489.490 1766.910 2490.670 ;
        RECT 1764.130 2311.090 1765.310 2312.270 ;
        RECT 1765.730 2311.090 1766.910 2312.270 ;
        RECT 1764.130 2309.490 1765.310 2310.670 ;
        RECT 1765.730 2309.490 1766.910 2310.670 ;
        RECT 1764.130 2131.090 1765.310 2132.270 ;
        RECT 1765.730 2131.090 1766.910 2132.270 ;
        RECT 1764.130 2129.490 1765.310 2130.670 ;
        RECT 1765.730 2129.490 1766.910 2130.670 ;
        RECT 1764.130 1951.090 1765.310 1952.270 ;
        RECT 1765.730 1951.090 1766.910 1952.270 ;
        RECT 1764.130 1949.490 1765.310 1950.670 ;
        RECT 1765.730 1949.490 1766.910 1950.670 ;
        RECT 1764.130 1771.090 1765.310 1772.270 ;
        RECT 1765.730 1771.090 1766.910 1772.270 ;
        RECT 1764.130 1769.490 1765.310 1770.670 ;
        RECT 1765.730 1769.490 1766.910 1770.670 ;
        RECT 1764.130 1591.090 1765.310 1592.270 ;
        RECT 1765.730 1591.090 1766.910 1592.270 ;
        RECT 1764.130 1589.490 1765.310 1590.670 ;
        RECT 1765.730 1589.490 1766.910 1590.670 ;
        RECT 1764.130 1411.090 1765.310 1412.270 ;
        RECT 1765.730 1411.090 1766.910 1412.270 ;
        RECT 1764.130 1409.490 1765.310 1410.670 ;
        RECT 1765.730 1409.490 1766.910 1410.670 ;
        RECT 1764.130 1231.090 1765.310 1232.270 ;
        RECT 1765.730 1231.090 1766.910 1232.270 ;
        RECT 1764.130 1229.490 1765.310 1230.670 ;
        RECT 1765.730 1229.490 1766.910 1230.670 ;
        RECT 1764.130 1051.090 1765.310 1052.270 ;
        RECT 1765.730 1051.090 1766.910 1052.270 ;
        RECT 1764.130 1049.490 1765.310 1050.670 ;
        RECT 1765.730 1049.490 1766.910 1050.670 ;
        RECT 1764.130 871.090 1765.310 872.270 ;
        RECT 1765.730 871.090 1766.910 872.270 ;
        RECT 1764.130 869.490 1765.310 870.670 ;
        RECT 1765.730 869.490 1766.910 870.670 ;
        RECT 1764.130 691.090 1765.310 692.270 ;
        RECT 1765.730 691.090 1766.910 692.270 ;
        RECT 1764.130 689.490 1765.310 690.670 ;
        RECT 1765.730 689.490 1766.910 690.670 ;
        RECT 1764.130 511.090 1765.310 512.270 ;
        RECT 1765.730 511.090 1766.910 512.270 ;
        RECT 1764.130 509.490 1765.310 510.670 ;
        RECT 1765.730 509.490 1766.910 510.670 ;
        RECT 1764.130 331.090 1765.310 332.270 ;
        RECT 1765.730 331.090 1766.910 332.270 ;
        RECT 1764.130 329.490 1765.310 330.670 ;
        RECT 1765.730 329.490 1766.910 330.670 ;
        RECT 1764.130 151.090 1765.310 152.270 ;
        RECT 1765.730 151.090 1766.910 152.270 ;
        RECT 1764.130 149.490 1765.310 150.670 ;
        RECT 1765.730 149.490 1766.910 150.670 ;
        RECT 1764.130 -33.260 1765.310 -32.080 ;
        RECT 1765.730 -33.260 1766.910 -32.080 ;
        RECT 1764.130 -34.860 1765.310 -33.680 ;
        RECT 1765.730 -34.860 1766.910 -33.680 ;
        RECT 1944.130 3553.360 1945.310 3554.540 ;
        RECT 1945.730 3553.360 1946.910 3554.540 ;
        RECT 1944.130 3551.760 1945.310 3552.940 ;
        RECT 1945.730 3551.760 1946.910 3552.940 ;
        RECT 1944.130 3391.090 1945.310 3392.270 ;
        RECT 1945.730 3391.090 1946.910 3392.270 ;
        RECT 1944.130 3389.490 1945.310 3390.670 ;
        RECT 1945.730 3389.490 1946.910 3390.670 ;
        RECT 1944.130 3211.090 1945.310 3212.270 ;
        RECT 1945.730 3211.090 1946.910 3212.270 ;
        RECT 1944.130 3209.490 1945.310 3210.670 ;
        RECT 1945.730 3209.490 1946.910 3210.670 ;
        RECT 1944.130 3031.090 1945.310 3032.270 ;
        RECT 1945.730 3031.090 1946.910 3032.270 ;
        RECT 1944.130 3029.490 1945.310 3030.670 ;
        RECT 1945.730 3029.490 1946.910 3030.670 ;
        RECT 1944.130 2851.090 1945.310 2852.270 ;
        RECT 1945.730 2851.090 1946.910 2852.270 ;
        RECT 1944.130 2849.490 1945.310 2850.670 ;
        RECT 1945.730 2849.490 1946.910 2850.670 ;
        RECT 1944.130 2671.090 1945.310 2672.270 ;
        RECT 1945.730 2671.090 1946.910 2672.270 ;
        RECT 1944.130 2669.490 1945.310 2670.670 ;
        RECT 1945.730 2669.490 1946.910 2670.670 ;
        RECT 1944.130 2491.090 1945.310 2492.270 ;
        RECT 1945.730 2491.090 1946.910 2492.270 ;
        RECT 1944.130 2489.490 1945.310 2490.670 ;
        RECT 1945.730 2489.490 1946.910 2490.670 ;
        RECT 1944.130 2311.090 1945.310 2312.270 ;
        RECT 1945.730 2311.090 1946.910 2312.270 ;
        RECT 1944.130 2309.490 1945.310 2310.670 ;
        RECT 1945.730 2309.490 1946.910 2310.670 ;
        RECT 1944.130 2131.090 1945.310 2132.270 ;
        RECT 1945.730 2131.090 1946.910 2132.270 ;
        RECT 1944.130 2129.490 1945.310 2130.670 ;
        RECT 1945.730 2129.490 1946.910 2130.670 ;
        RECT 1944.130 1951.090 1945.310 1952.270 ;
        RECT 1945.730 1951.090 1946.910 1952.270 ;
        RECT 1944.130 1949.490 1945.310 1950.670 ;
        RECT 1945.730 1949.490 1946.910 1950.670 ;
        RECT 1944.130 1771.090 1945.310 1772.270 ;
        RECT 1945.730 1771.090 1946.910 1772.270 ;
        RECT 1944.130 1769.490 1945.310 1770.670 ;
        RECT 1945.730 1769.490 1946.910 1770.670 ;
        RECT 1944.130 1591.090 1945.310 1592.270 ;
        RECT 1945.730 1591.090 1946.910 1592.270 ;
        RECT 1944.130 1589.490 1945.310 1590.670 ;
        RECT 1945.730 1589.490 1946.910 1590.670 ;
        RECT 1944.130 1411.090 1945.310 1412.270 ;
        RECT 1945.730 1411.090 1946.910 1412.270 ;
        RECT 1944.130 1409.490 1945.310 1410.670 ;
        RECT 1945.730 1409.490 1946.910 1410.670 ;
        RECT 1944.130 1231.090 1945.310 1232.270 ;
        RECT 1945.730 1231.090 1946.910 1232.270 ;
        RECT 1944.130 1229.490 1945.310 1230.670 ;
        RECT 1945.730 1229.490 1946.910 1230.670 ;
        RECT 1944.130 1051.090 1945.310 1052.270 ;
        RECT 1945.730 1051.090 1946.910 1052.270 ;
        RECT 1944.130 1049.490 1945.310 1050.670 ;
        RECT 1945.730 1049.490 1946.910 1050.670 ;
        RECT 1944.130 871.090 1945.310 872.270 ;
        RECT 1945.730 871.090 1946.910 872.270 ;
        RECT 1944.130 869.490 1945.310 870.670 ;
        RECT 1945.730 869.490 1946.910 870.670 ;
        RECT 1944.130 691.090 1945.310 692.270 ;
        RECT 1945.730 691.090 1946.910 692.270 ;
        RECT 1944.130 689.490 1945.310 690.670 ;
        RECT 1945.730 689.490 1946.910 690.670 ;
        RECT 1944.130 511.090 1945.310 512.270 ;
        RECT 1945.730 511.090 1946.910 512.270 ;
        RECT 1944.130 509.490 1945.310 510.670 ;
        RECT 1945.730 509.490 1946.910 510.670 ;
        RECT 1944.130 331.090 1945.310 332.270 ;
        RECT 1945.730 331.090 1946.910 332.270 ;
        RECT 1944.130 329.490 1945.310 330.670 ;
        RECT 1945.730 329.490 1946.910 330.670 ;
        RECT 1944.130 151.090 1945.310 152.270 ;
        RECT 1945.730 151.090 1946.910 152.270 ;
        RECT 1944.130 149.490 1945.310 150.670 ;
        RECT 1945.730 149.490 1946.910 150.670 ;
        RECT 1944.130 -33.260 1945.310 -32.080 ;
        RECT 1945.730 -33.260 1946.910 -32.080 ;
        RECT 1944.130 -34.860 1945.310 -33.680 ;
        RECT 1945.730 -34.860 1946.910 -33.680 ;
        RECT 2124.130 3553.360 2125.310 3554.540 ;
        RECT 2125.730 3553.360 2126.910 3554.540 ;
        RECT 2124.130 3551.760 2125.310 3552.940 ;
        RECT 2125.730 3551.760 2126.910 3552.940 ;
        RECT 2124.130 3391.090 2125.310 3392.270 ;
        RECT 2125.730 3391.090 2126.910 3392.270 ;
        RECT 2124.130 3389.490 2125.310 3390.670 ;
        RECT 2125.730 3389.490 2126.910 3390.670 ;
        RECT 2124.130 3211.090 2125.310 3212.270 ;
        RECT 2125.730 3211.090 2126.910 3212.270 ;
        RECT 2124.130 3209.490 2125.310 3210.670 ;
        RECT 2125.730 3209.490 2126.910 3210.670 ;
        RECT 2124.130 3031.090 2125.310 3032.270 ;
        RECT 2125.730 3031.090 2126.910 3032.270 ;
        RECT 2124.130 3029.490 2125.310 3030.670 ;
        RECT 2125.730 3029.490 2126.910 3030.670 ;
        RECT 2124.130 2851.090 2125.310 2852.270 ;
        RECT 2125.730 2851.090 2126.910 2852.270 ;
        RECT 2124.130 2849.490 2125.310 2850.670 ;
        RECT 2125.730 2849.490 2126.910 2850.670 ;
        RECT 2124.130 2671.090 2125.310 2672.270 ;
        RECT 2125.730 2671.090 2126.910 2672.270 ;
        RECT 2124.130 2669.490 2125.310 2670.670 ;
        RECT 2125.730 2669.490 2126.910 2670.670 ;
        RECT 2124.130 2491.090 2125.310 2492.270 ;
        RECT 2125.730 2491.090 2126.910 2492.270 ;
        RECT 2124.130 2489.490 2125.310 2490.670 ;
        RECT 2125.730 2489.490 2126.910 2490.670 ;
        RECT 2124.130 2311.090 2125.310 2312.270 ;
        RECT 2125.730 2311.090 2126.910 2312.270 ;
        RECT 2124.130 2309.490 2125.310 2310.670 ;
        RECT 2125.730 2309.490 2126.910 2310.670 ;
        RECT 2124.130 2131.090 2125.310 2132.270 ;
        RECT 2125.730 2131.090 2126.910 2132.270 ;
        RECT 2124.130 2129.490 2125.310 2130.670 ;
        RECT 2125.730 2129.490 2126.910 2130.670 ;
        RECT 2124.130 1951.090 2125.310 1952.270 ;
        RECT 2125.730 1951.090 2126.910 1952.270 ;
        RECT 2124.130 1949.490 2125.310 1950.670 ;
        RECT 2125.730 1949.490 2126.910 1950.670 ;
        RECT 2124.130 1771.090 2125.310 1772.270 ;
        RECT 2125.730 1771.090 2126.910 1772.270 ;
        RECT 2124.130 1769.490 2125.310 1770.670 ;
        RECT 2125.730 1769.490 2126.910 1770.670 ;
        RECT 2124.130 1591.090 2125.310 1592.270 ;
        RECT 2125.730 1591.090 2126.910 1592.270 ;
        RECT 2124.130 1589.490 2125.310 1590.670 ;
        RECT 2125.730 1589.490 2126.910 1590.670 ;
        RECT 2124.130 1411.090 2125.310 1412.270 ;
        RECT 2125.730 1411.090 2126.910 1412.270 ;
        RECT 2124.130 1409.490 2125.310 1410.670 ;
        RECT 2125.730 1409.490 2126.910 1410.670 ;
        RECT 2124.130 1231.090 2125.310 1232.270 ;
        RECT 2125.730 1231.090 2126.910 1232.270 ;
        RECT 2124.130 1229.490 2125.310 1230.670 ;
        RECT 2125.730 1229.490 2126.910 1230.670 ;
        RECT 2124.130 1051.090 2125.310 1052.270 ;
        RECT 2125.730 1051.090 2126.910 1052.270 ;
        RECT 2124.130 1049.490 2125.310 1050.670 ;
        RECT 2125.730 1049.490 2126.910 1050.670 ;
        RECT 2124.130 871.090 2125.310 872.270 ;
        RECT 2125.730 871.090 2126.910 872.270 ;
        RECT 2124.130 869.490 2125.310 870.670 ;
        RECT 2125.730 869.490 2126.910 870.670 ;
        RECT 2124.130 691.090 2125.310 692.270 ;
        RECT 2125.730 691.090 2126.910 692.270 ;
        RECT 2124.130 689.490 2125.310 690.670 ;
        RECT 2125.730 689.490 2126.910 690.670 ;
        RECT 2124.130 511.090 2125.310 512.270 ;
        RECT 2125.730 511.090 2126.910 512.270 ;
        RECT 2124.130 509.490 2125.310 510.670 ;
        RECT 2125.730 509.490 2126.910 510.670 ;
        RECT 2124.130 331.090 2125.310 332.270 ;
        RECT 2125.730 331.090 2126.910 332.270 ;
        RECT 2124.130 329.490 2125.310 330.670 ;
        RECT 2125.730 329.490 2126.910 330.670 ;
        RECT 2124.130 151.090 2125.310 152.270 ;
        RECT 2125.730 151.090 2126.910 152.270 ;
        RECT 2124.130 149.490 2125.310 150.670 ;
        RECT 2125.730 149.490 2126.910 150.670 ;
        RECT 2124.130 -33.260 2125.310 -32.080 ;
        RECT 2125.730 -33.260 2126.910 -32.080 ;
        RECT 2124.130 -34.860 2125.310 -33.680 ;
        RECT 2125.730 -34.860 2126.910 -33.680 ;
        RECT 2304.130 3553.360 2305.310 3554.540 ;
        RECT 2305.730 3553.360 2306.910 3554.540 ;
        RECT 2304.130 3551.760 2305.310 3552.940 ;
        RECT 2305.730 3551.760 2306.910 3552.940 ;
        RECT 2304.130 3391.090 2305.310 3392.270 ;
        RECT 2305.730 3391.090 2306.910 3392.270 ;
        RECT 2304.130 3389.490 2305.310 3390.670 ;
        RECT 2305.730 3389.490 2306.910 3390.670 ;
        RECT 2304.130 3211.090 2305.310 3212.270 ;
        RECT 2305.730 3211.090 2306.910 3212.270 ;
        RECT 2304.130 3209.490 2305.310 3210.670 ;
        RECT 2305.730 3209.490 2306.910 3210.670 ;
        RECT 2304.130 3031.090 2305.310 3032.270 ;
        RECT 2305.730 3031.090 2306.910 3032.270 ;
        RECT 2304.130 3029.490 2305.310 3030.670 ;
        RECT 2305.730 3029.490 2306.910 3030.670 ;
        RECT 2304.130 2851.090 2305.310 2852.270 ;
        RECT 2305.730 2851.090 2306.910 2852.270 ;
        RECT 2304.130 2849.490 2305.310 2850.670 ;
        RECT 2305.730 2849.490 2306.910 2850.670 ;
        RECT 2304.130 2671.090 2305.310 2672.270 ;
        RECT 2305.730 2671.090 2306.910 2672.270 ;
        RECT 2304.130 2669.490 2305.310 2670.670 ;
        RECT 2305.730 2669.490 2306.910 2670.670 ;
        RECT 2304.130 2491.090 2305.310 2492.270 ;
        RECT 2305.730 2491.090 2306.910 2492.270 ;
        RECT 2304.130 2489.490 2305.310 2490.670 ;
        RECT 2305.730 2489.490 2306.910 2490.670 ;
        RECT 2304.130 2311.090 2305.310 2312.270 ;
        RECT 2305.730 2311.090 2306.910 2312.270 ;
        RECT 2304.130 2309.490 2305.310 2310.670 ;
        RECT 2305.730 2309.490 2306.910 2310.670 ;
        RECT 2304.130 2131.090 2305.310 2132.270 ;
        RECT 2305.730 2131.090 2306.910 2132.270 ;
        RECT 2304.130 2129.490 2305.310 2130.670 ;
        RECT 2305.730 2129.490 2306.910 2130.670 ;
        RECT 2304.130 1951.090 2305.310 1952.270 ;
        RECT 2305.730 1951.090 2306.910 1952.270 ;
        RECT 2304.130 1949.490 2305.310 1950.670 ;
        RECT 2305.730 1949.490 2306.910 1950.670 ;
        RECT 2304.130 1771.090 2305.310 1772.270 ;
        RECT 2305.730 1771.090 2306.910 1772.270 ;
        RECT 2304.130 1769.490 2305.310 1770.670 ;
        RECT 2305.730 1769.490 2306.910 1770.670 ;
        RECT 2304.130 1591.090 2305.310 1592.270 ;
        RECT 2305.730 1591.090 2306.910 1592.270 ;
        RECT 2304.130 1589.490 2305.310 1590.670 ;
        RECT 2305.730 1589.490 2306.910 1590.670 ;
        RECT 2304.130 1411.090 2305.310 1412.270 ;
        RECT 2305.730 1411.090 2306.910 1412.270 ;
        RECT 2304.130 1409.490 2305.310 1410.670 ;
        RECT 2305.730 1409.490 2306.910 1410.670 ;
        RECT 2304.130 1231.090 2305.310 1232.270 ;
        RECT 2305.730 1231.090 2306.910 1232.270 ;
        RECT 2304.130 1229.490 2305.310 1230.670 ;
        RECT 2305.730 1229.490 2306.910 1230.670 ;
        RECT 2304.130 1051.090 2305.310 1052.270 ;
        RECT 2305.730 1051.090 2306.910 1052.270 ;
        RECT 2304.130 1049.490 2305.310 1050.670 ;
        RECT 2305.730 1049.490 2306.910 1050.670 ;
        RECT 2304.130 871.090 2305.310 872.270 ;
        RECT 2305.730 871.090 2306.910 872.270 ;
        RECT 2304.130 869.490 2305.310 870.670 ;
        RECT 2305.730 869.490 2306.910 870.670 ;
        RECT 2304.130 691.090 2305.310 692.270 ;
        RECT 2305.730 691.090 2306.910 692.270 ;
        RECT 2304.130 689.490 2305.310 690.670 ;
        RECT 2305.730 689.490 2306.910 690.670 ;
        RECT 2304.130 511.090 2305.310 512.270 ;
        RECT 2305.730 511.090 2306.910 512.270 ;
        RECT 2304.130 509.490 2305.310 510.670 ;
        RECT 2305.730 509.490 2306.910 510.670 ;
        RECT 2304.130 331.090 2305.310 332.270 ;
        RECT 2305.730 331.090 2306.910 332.270 ;
        RECT 2304.130 329.490 2305.310 330.670 ;
        RECT 2305.730 329.490 2306.910 330.670 ;
        RECT 2304.130 151.090 2305.310 152.270 ;
        RECT 2305.730 151.090 2306.910 152.270 ;
        RECT 2304.130 149.490 2305.310 150.670 ;
        RECT 2305.730 149.490 2306.910 150.670 ;
        RECT 2304.130 -33.260 2305.310 -32.080 ;
        RECT 2305.730 -33.260 2306.910 -32.080 ;
        RECT 2304.130 -34.860 2305.310 -33.680 ;
        RECT 2305.730 -34.860 2306.910 -33.680 ;
        RECT 2484.130 3553.360 2485.310 3554.540 ;
        RECT 2485.730 3553.360 2486.910 3554.540 ;
        RECT 2484.130 3551.760 2485.310 3552.940 ;
        RECT 2485.730 3551.760 2486.910 3552.940 ;
        RECT 2484.130 3391.090 2485.310 3392.270 ;
        RECT 2485.730 3391.090 2486.910 3392.270 ;
        RECT 2484.130 3389.490 2485.310 3390.670 ;
        RECT 2485.730 3389.490 2486.910 3390.670 ;
        RECT 2484.130 3211.090 2485.310 3212.270 ;
        RECT 2485.730 3211.090 2486.910 3212.270 ;
        RECT 2484.130 3209.490 2485.310 3210.670 ;
        RECT 2485.730 3209.490 2486.910 3210.670 ;
        RECT 2484.130 3031.090 2485.310 3032.270 ;
        RECT 2485.730 3031.090 2486.910 3032.270 ;
        RECT 2484.130 3029.490 2485.310 3030.670 ;
        RECT 2485.730 3029.490 2486.910 3030.670 ;
        RECT 2484.130 2851.090 2485.310 2852.270 ;
        RECT 2485.730 2851.090 2486.910 2852.270 ;
        RECT 2484.130 2849.490 2485.310 2850.670 ;
        RECT 2485.730 2849.490 2486.910 2850.670 ;
        RECT 2484.130 2671.090 2485.310 2672.270 ;
        RECT 2485.730 2671.090 2486.910 2672.270 ;
        RECT 2484.130 2669.490 2485.310 2670.670 ;
        RECT 2485.730 2669.490 2486.910 2670.670 ;
        RECT 2484.130 2491.090 2485.310 2492.270 ;
        RECT 2485.730 2491.090 2486.910 2492.270 ;
        RECT 2484.130 2489.490 2485.310 2490.670 ;
        RECT 2485.730 2489.490 2486.910 2490.670 ;
        RECT 2484.130 2311.090 2485.310 2312.270 ;
        RECT 2485.730 2311.090 2486.910 2312.270 ;
        RECT 2484.130 2309.490 2485.310 2310.670 ;
        RECT 2485.730 2309.490 2486.910 2310.670 ;
        RECT 2484.130 2131.090 2485.310 2132.270 ;
        RECT 2485.730 2131.090 2486.910 2132.270 ;
        RECT 2484.130 2129.490 2485.310 2130.670 ;
        RECT 2485.730 2129.490 2486.910 2130.670 ;
        RECT 2484.130 1951.090 2485.310 1952.270 ;
        RECT 2485.730 1951.090 2486.910 1952.270 ;
        RECT 2484.130 1949.490 2485.310 1950.670 ;
        RECT 2485.730 1949.490 2486.910 1950.670 ;
        RECT 2484.130 1771.090 2485.310 1772.270 ;
        RECT 2485.730 1771.090 2486.910 1772.270 ;
        RECT 2484.130 1769.490 2485.310 1770.670 ;
        RECT 2485.730 1769.490 2486.910 1770.670 ;
        RECT 2484.130 1591.090 2485.310 1592.270 ;
        RECT 2485.730 1591.090 2486.910 1592.270 ;
        RECT 2484.130 1589.490 2485.310 1590.670 ;
        RECT 2485.730 1589.490 2486.910 1590.670 ;
        RECT 2484.130 1411.090 2485.310 1412.270 ;
        RECT 2485.730 1411.090 2486.910 1412.270 ;
        RECT 2484.130 1409.490 2485.310 1410.670 ;
        RECT 2485.730 1409.490 2486.910 1410.670 ;
        RECT 2484.130 1231.090 2485.310 1232.270 ;
        RECT 2485.730 1231.090 2486.910 1232.270 ;
        RECT 2484.130 1229.490 2485.310 1230.670 ;
        RECT 2485.730 1229.490 2486.910 1230.670 ;
        RECT 2484.130 1051.090 2485.310 1052.270 ;
        RECT 2485.730 1051.090 2486.910 1052.270 ;
        RECT 2484.130 1049.490 2485.310 1050.670 ;
        RECT 2485.730 1049.490 2486.910 1050.670 ;
        RECT 2484.130 871.090 2485.310 872.270 ;
        RECT 2485.730 871.090 2486.910 872.270 ;
        RECT 2484.130 869.490 2485.310 870.670 ;
        RECT 2485.730 869.490 2486.910 870.670 ;
        RECT 2484.130 691.090 2485.310 692.270 ;
        RECT 2485.730 691.090 2486.910 692.270 ;
        RECT 2484.130 689.490 2485.310 690.670 ;
        RECT 2485.730 689.490 2486.910 690.670 ;
        RECT 2484.130 511.090 2485.310 512.270 ;
        RECT 2485.730 511.090 2486.910 512.270 ;
        RECT 2484.130 509.490 2485.310 510.670 ;
        RECT 2485.730 509.490 2486.910 510.670 ;
        RECT 2484.130 331.090 2485.310 332.270 ;
        RECT 2485.730 331.090 2486.910 332.270 ;
        RECT 2484.130 329.490 2485.310 330.670 ;
        RECT 2485.730 329.490 2486.910 330.670 ;
        RECT 2484.130 151.090 2485.310 152.270 ;
        RECT 2485.730 151.090 2486.910 152.270 ;
        RECT 2484.130 149.490 2485.310 150.670 ;
        RECT 2485.730 149.490 2486.910 150.670 ;
        RECT 2484.130 -33.260 2485.310 -32.080 ;
        RECT 2485.730 -33.260 2486.910 -32.080 ;
        RECT 2484.130 -34.860 2485.310 -33.680 ;
        RECT 2485.730 -34.860 2486.910 -33.680 ;
        RECT 2664.130 3553.360 2665.310 3554.540 ;
        RECT 2665.730 3553.360 2666.910 3554.540 ;
        RECT 2664.130 3551.760 2665.310 3552.940 ;
        RECT 2665.730 3551.760 2666.910 3552.940 ;
        RECT 2664.130 3391.090 2665.310 3392.270 ;
        RECT 2665.730 3391.090 2666.910 3392.270 ;
        RECT 2664.130 3389.490 2665.310 3390.670 ;
        RECT 2665.730 3389.490 2666.910 3390.670 ;
        RECT 2664.130 3211.090 2665.310 3212.270 ;
        RECT 2665.730 3211.090 2666.910 3212.270 ;
        RECT 2664.130 3209.490 2665.310 3210.670 ;
        RECT 2665.730 3209.490 2666.910 3210.670 ;
        RECT 2664.130 3031.090 2665.310 3032.270 ;
        RECT 2665.730 3031.090 2666.910 3032.270 ;
        RECT 2664.130 3029.490 2665.310 3030.670 ;
        RECT 2665.730 3029.490 2666.910 3030.670 ;
        RECT 2664.130 2851.090 2665.310 2852.270 ;
        RECT 2665.730 2851.090 2666.910 2852.270 ;
        RECT 2664.130 2849.490 2665.310 2850.670 ;
        RECT 2665.730 2849.490 2666.910 2850.670 ;
        RECT 2664.130 2671.090 2665.310 2672.270 ;
        RECT 2665.730 2671.090 2666.910 2672.270 ;
        RECT 2664.130 2669.490 2665.310 2670.670 ;
        RECT 2665.730 2669.490 2666.910 2670.670 ;
        RECT 2664.130 2491.090 2665.310 2492.270 ;
        RECT 2665.730 2491.090 2666.910 2492.270 ;
        RECT 2664.130 2489.490 2665.310 2490.670 ;
        RECT 2665.730 2489.490 2666.910 2490.670 ;
        RECT 2664.130 2311.090 2665.310 2312.270 ;
        RECT 2665.730 2311.090 2666.910 2312.270 ;
        RECT 2664.130 2309.490 2665.310 2310.670 ;
        RECT 2665.730 2309.490 2666.910 2310.670 ;
        RECT 2664.130 2131.090 2665.310 2132.270 ;
        RECT 2665.730 2131.090 2666.910 2132.270 ;
        RECT 2664.130 2129.490 2665.310 2130.670 ;
        RECT 2665.730 2129.490 2666.910 2130.670 ;
        RECT 2664.130 1951.090 2665.310 1952.270 ;
        RECT 2665.730 1951.090 2666.910 1952.270 ;
        RECT 2664.130 1949.490 2665.310 1950.670 ;
        RECT 2665.730 1949.490 2666.910 1950.670 ;
        RECT 2664.130 1771.090 2665.310 1772.270 ;
        RECT 2665.730 1771.090 2666.910 1772.270 ;
        RECT 2664.130 1769.490 2665.310 1770.670 ;
        RECT 2665.730 1769.490 2666.910 1770.670 ;
        RECT 2664.130 1591.090 2665.310 1592.270 ;
        RECT 2665.730 1591.090 2666.910 1592.270 ;
        RECT 2664.130 1589.490 2665.310 1590.670 ;
        RECT 2665.730 1589.490 2666.910 1590.670 ;
        RECT 2664.130 1411.090 2665.310 1412.270 ;
        RECT 2665.730 1411.090 2666.910 1412.270 ;
        RECT 2664.130 1409.490 2665.310 1410.670 ;
        RECT 2665.730 1409.490 2666.910 1410.670 ;
        RECT 2664.130 1231.090 2665.310 1232.270 ;
        RECT 2665.730 1231.090 2666.910 1232.270 ;
        RECT 2664.130 1229.490 2665.310 1230.670 ;
        RECT 2665.730 1229.490 2666.910 1230.670 ;
        RECT 2664.130 1051.090 2665.310 1052.270 ;
        RECT 2665.730 1051.090 2666.910 1052.270 ;
        RECT 2664.130 1049.490 2665.310 1050.670 ;
        RECT 2665.730 1049.490 2666.910 1050.670 ;
        RECT 2664.130 871.090 2665.310 872.270 ;
        RECT 2665.730 871.090 2666.910 872.270 ;
        RECT 2664.130 869.490 2665.310 870.670 ;
        RECT 2665.730 869.490 2666.910 870.670 ;
        RECT 2664.130 691.090 2665.310 692.270 ;
        RECT 2665.730 691.090 2666.910 692.270 ;
        RECT 2664.130 689.490 2665.310 690.670 ;
        RECT 2665.730 689.490 2666.910 690.670 ;
        RECT 2664.130 511.090 2665.310 512.270 ;
        RECT 2665.730 511.090 2666.910 512.270 ;
        RECT 2664.130 509.490 2665.310 510.670 ;
        RECT 2665.730 509.490 2666.910 510.670 ;
        RECT 2664.130 331.090 2665.310 332.270 ;
        RECT 2665.730 331.090 2666.910 332.270 ;
        RECT 2664.130 329.490 2665.310 330.670 ;
        RECT 2665.730 329.490 2666.910 330.670 ;
        RECT 2664.130 151.090 2665.310 152.270 ;
        RECT 2665.730 151.090 2666.910 152.270 ;
        RECT 2664.130 149.490 2665.310 150.670 ;
        RECT 2665.730 149.490 2666.910 150.670 ;
        RECT 2664.130 -33.260 2665.310 -32.080 ;
        RECT 2665.730 -33.260 2666.910 -32.080 ;
        RECT 2664.130 -34.860 2665.310 -33.680 ;
        RECT 2665.730 -34.860 2666.910 -33.680 ;
        RECT 2844.130 3553.360 2845.310 3554.540 ;
        RECT 2845.730 3553.360 2846.910 3554.540 ;
        RECT 2844.130 3551.760 2845.310 3552.940 ;
        RECT 2845.730 3551.760 2846.910 3552.940 ;
        RECT 2844.130 3391.090 2845.310 3392.270 ;
        RECT 2845.730 3391.090 2846.910 3392.270 ;
        RECT 2844.130 3389.490 2845.310 3390.670 ;
        RECT 2845.730 3389.490 2846.910 3390.670 ;
        RECT 2844.130 3211.090 2845.310 3212.270 ;
        RECT 2845.730 3211.090 2846.910 3212.270 ;
        RECT 2844.130 3209.490 2845.310 3210.670 ;
        RECT 2845.730 3209.490 2846.910 3210.670 ;
        RECT 2844.130 3031.090 2845.310 3032.270 ;
        RECT 2845.730 3031.090 2846.910 3032.270 ;
        RECT 2844.130 3029.490 2845.310 3030.670 ;
        RECT 2845.730 3029.490 2846.910 3030.670 ;
        RECT 2844.130 2851.090 2845.310 2852.270 ;
        RECT 2845.730 2851.090 2846.910 2852.270 ;
        RECT 2844.130 2849.490 2845.310 2850.670 ;
        RECT 2845.730 2849.490 2846.910 2850.670 ;
        RECT 2844.130 2671.090 2845.310 2672.270 ;
        RECT 2845.730 2671.090 2846.910 2672.270 ;
        RECT 2844.130 2669.490 2845.310 2670.670 ;
        RECT 2845.730 2669.490 2846.910 2670.670 ;
        RECT 2844.130 2491.090 2845.310 2492.270 ;
        RECT 2845.730 2491.090 2846.910 2492.270 ;
        RECT 2844.130 2489.490 2845.310 2490.670 ;
        RECT 2845.730 2489.490 2846.910 2490.670 ;
        RECT 2844.130 2311.090 2845.310 2312.270 ;
        RECT 2845.730 2311.090 2846.910 2312.270 ;
        RECT 2844.130 2309.490 2845.310 2310.670 ;
        RECT 2845.730 2309.490 2846.910 2310.670 ;
        RECT 2844.130 2131.090 2845.310 2132.270 ;
        RECT 2845.730 2131.090 2846.910 2132.270 ;
        RECT 2844.130 2129.490 2845.310 2130.670 ;
        RECT 2845.730 2129.490 2846.910 2130.670 ;
        RECT 2844.130 1951.090 2845.310 1952.270 ;
        RECT 2845.730 1951.090 2846.910 1952.270 ;
        RECT 2844.130 1949.490 2845.310 1950.670 ;
        RECT 2845.730 1949.490 2846.910 1950.670 ;
        RECT 2844.130 1771.090 2845.310 1772.270 ;
        RECT 2845.730 1771.090 2846.910 1772.270 ;
        RECT 2844.130 1769.490 2845.310 1770.670 ;
        RECT 2845.730 1769.490 2846.910 1770.670 ;
        RECT 2844.130 1591.090 2845.310 1592.270 ;
        RECT 2845.730 1591.090 2846.910 1592.270 ;
        RECT 2844.130 1589.490 2845.310 1590.670 ;
        RECT 2845.730 1589.490 2846.910 1590.670 ;
        RECT 2844.130 1411.090 2845.310 1412.270 ;
        RECT 2845.730 1411.090 2846.910 1412.270 ;
        RECT 2844.130 1409.490 2845.310 1410.670 ;
        RECT 2845.730 1409.490 2846.910 1410.670 ;
        RECT 2844.130 1231.090 2845.310 1232.270 ;
        RECT 2845.730 1231.090 2846.910 1232.270 ;
        RECT 2844.130 1229.490 2845.310 1230.670 ;
        RECT 2845.730 1229.490 2846.910 1230.670 ;
        RECT 2844.130 1051.090 2845.310 1052.270 ;
        RECT 2845.730 1051.090 2846.910 1052.270 ;
        RECT 2844.130 1049.490 2845.310 1050.670 ;
        RECT 2845.730 1049.490 2846.910 1050.670 ;
        RECT 2844.130 871.090 2845.310 872.270 ;
        RECT 2845.730 871.090 2846.910 872.270 ;
        RECT 2844.130 869.490 2845.310 870.670 ;
        RECT 2845.730 869.490 2846.910 870.670 ;
        RECT 2844.130 691.090 2845.310 692.270 ;
        RECT 2845.730 691.090 2846.910 692.270 ;
        RECT 2844.130 689.490 2845.310 690.670 ;
        RECT 2845.730 689.490 2846.910 690.670 ;
        RECT 2844.130 511.090 2845.310 512.270 ;
        RECT 2845.730 511.090 2846.910 512.270 ;
        RECT 2844.130 509.490 2845.310 510.670 ;
        RECT 2845.730 509.490 2846.910 510.670 ;
        RECT 2844.130 331.090 2845.310 332.270 ;
        RECT 2845.730 331.090 2846.910 332.270 ;
        RECT 2844.130 329.490 2845.310 330.670 ;
        RECT 2845.730 329.490 2846.910 330.670 ;
        RECT 2844.130 151.090 2845.310 152.270 ;
        RECT 2845.730 151.090 2846.910 152.270 ;
        RECT 2844.130 149.490 2845.310 150.670 ;
        RECT 2845.730 149.490 2846.910 150.670 ;
        RECT 2844.130 -33.260 2845.310 -32.080 ;
        RECT 2845.730 -33.260 2846.910 -32.080 ;
        RECT 2844.130 -34.860 2845.310 -33.680 ;
        RECT 2845.730 -34.860 2846.910 -33.680 ;
        RECT 2957.060 3553.360 2958.240 3554.540 ;
        RECT 2958.660 3553.360 2959.840 3554.540 ;
        RECT 2957.060 3551.760 2958.240 3552.940 ;
        RECT 2958.660 3551.760 2959.840 3552.940 ;
        RECT 2957.060 3391.090 2958.240 3392.270 ;
        RECT 2958.660 3391.090 2959.840 3392.270 ;
        RECT 2957.060 3389.490 2958.240 3390.670 ;
        RECT 2958.660 3389.490 2959.840 3390.670 ;
        RECT 2957.060 3211.090 2958.240 3212.270 ;
        RECT 2958.660 3211.090 2959.840 3212.270 ;
        RECT 2957.060 3209.490 2958.240 3210.670 ;
        RECT 2958.660 3209.490 2959.840 3210.670 ;
        RECT 2957.060 3031.090 2958.240 3032.270 ;
        RECT 2958.660 3031.090 2959.840 3032.270 ;
        RECT 2957.060 3029.490 2958.240 3030.670 ;
        RECT 2958.660 3029.490 2959.840 3030.670 ;
        RECT 2957.060 2851.090 2958.240 2852.270 ;
        RECT 2958.660 2851.090 2959.840 2852.270 ;
        RECT 2957.060 2849.490 2958.240 2850.670 ;
        RECT 2958.660 2849.490 2959.840 2850.670 ;
        RECT 2957.060 2671.090 2958.240 2672.270 ;
        RECT 2958.660 2671.090 2959.840 2672.270 ;
        RECT 2957.060 2669.490 2958.240 2670.670 ;
        RECT 2958.660 2669.490 2959.840 2670.670 ;
        RECT 2957.060 2491.090 2958.240 2492.270 ;
        RECT 2958.660 2491.090 2959.840 2492.270 ;
        RECT 2957.060 2489.490 2958.240 2490.670 ;
        RECT 2958.660 2489.490 2959.840 2490.670 ;
        RECT 2957.060 2311.090 2958.240 2312.270 ;
        RECT 2958.660 2311.090 2959.840 2312.270 ;
        RECT 2957.060 2309.490 2958.240 2310.670 ;
        RECT 2958.660 2309.490 2959.840 2310.670 ;
        RECT 2957.060 2131.090 2958.240 2132.270 ;
        RECT 2958.660 2131.090 2959.840 2132.270 ;
        RECT 2957.060 2129.490 2958.240 2130.670 ;
        RECT 2958.660 2129.490 2959.840 2130.670 ;
        RECT 2957.060 1951.090 2958.240 1952.270 ;
        RECT 2958.660 1951.090 2959.840 1952.270 ;
        RECT 2957.060 1949.490 2958.240 1950.670 ;
        RECT 2958.660 1949.490 2959.840 1950.670 ;
        RECT 2957.060 1771.090 2958.240 1772.270 ;
        RECT 2958.660 1771.090 2959.840 1772.270 ;
        RECT 2957.060 1769.490 2958.240 1770.670 ;
        RECT 2958.660 1769.490 2959.840 1770.670 ;
        RECT 2957.060 1591.090 2958.240 1592.270 ;
        RECT 2958.660 1591.090 2959.840 1592.270 ;
        RECT 2957.060 1589.490 2958.240 1590.670 ;
        RECT 2958.660 1589.490 2959.840 1590.670 ;
        RECT 2957.060 1411.090 2958.240 1412.270 ;
        RECT 2958.660 1411.090 2959.840 1412.270 ;
        RECT 2957.060 1409.490 2958.240 1410.670 ;
        RECT 2958.660 1409.490 2959.840 1410.670 ;
        RECT 2957.060 1231.090 2958.240 1232.270 ;
        RECT 2958.660 1231.090 2959.840 1232.270 ;
        RECT 2957.060 1229.490 2958.240 1230.670 ;
        RECT 2958.660 1229.490 2959.840 1230.670 ;
        RECT 2957.060 1051.090 2958.240 1052.270 ;
        RECT 2958.660 1051.090 2959.840 1052.270 ;
        RECT 2957.060 1049.490 2958.240 1050.670 ;
        RECT 2958.660 1049.490 2959.840 1050.670 ;
        RECT 2957.060 871.090 2958.240 872.270 ;
        RECT 2958.660 871.090 2959.840 872.270 ;
        RECT 2957.060 869.490 2958.240 870.670 ;
        RECT 2958.660 869.490 2959.840 870.670 ;
        RECT 2957.060 691.090 2958.240 692.270 ;
        RECT 2958.660 691.090 2959.840 692.270 ;
        RECT 2957.060 689.490 2958.240 690.670 ;
        RECT 2958.660 689.490 2959.840 690.670 ;
        RECT 2957.060 511.090 2958.240 512.270 ;
        RECT 2958.660 511.090 2959.840 512.270 ;
        RECT 2957.060 509.490 2958.240 510.670 ;
        RECT 2958.660 509.490 2959.840 510.670 ;
        RECT 2957.060 331.090 2958.240 332.270 ;
        RECT 2958.660 331.090 2959.840 332.270 ;
        RECT 2957.060 329.490 2958.240 330.670 ;
        RECT 2958.660 329.490 2959.840 330.670 ;
        RECT 2957.060 151.090 2958.240 152.270 ;
        RECT 2958.660 151.090 2959.840 152.270 ;
        RECT 2957.060 149.490 2958.240 150.670 ;
        RECT 2958.660 149.490 2959.840 150.670 ;
        RECT 2957.060 -33.260 2958.240 -32.080 ;
        RECT 2958.660 -33.260 2959.840 -32.080 ;
        RECT 2957.060 -34.860 2958.240 -33.680 ;
        RECT 2958.660 -34.860 2959.840 -33.680 ;
      LAYER met5 ;
        RECT -40.380 3551.600 2960.000 3554.700 ;
        RECT -45.180 3389.330 2964.800 3392.430 ;
        RECT -45.180 3209.330 2964.800 3212.430 ;
        RECT -45.180 3029.330 2964.800 3032.430 ;
        RECT -45.180 2849.330 2964.800 2852.430 ;
        RECT -45.180 2669.330 2964.800 2672.430 ;
        RECT -45.180 2489.330 2964.800 2492.430 ;
        RECT -45.180 2309.330 2964.800 2312.430 ;
        RECT -45.180 2129.330 2964.800 2132.430 ;
        RECT -45.180 1949.330 2964.800 1952.430 ;
        RECT -45.180 1769.330 2964.800 1772.430 ;
        RECT -45.180 1589.330 2964.800 1592.430 ;
        RECT -45.180 1409.330 2964.800 1412.430 ;
        RECT -45.180 1229.330 2964.800 1232.430 ;
        RECT -45.180 1049.330 2964.800 1052.430 ;
        RECT -45.180 869.330 2964.800 872.430 ;
        RECT -45.180 689.330 2964.800 692.430 ;
        RECT -45.180 509.330 2964.800 512.430 ;
        RECT -45.180 329.330 2964.800 332.430 ;
        RECT -45.180 149.330 2964.800 152.430 ;
        RECT -40.380 -35.020 2960.000 -31.920 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -35.580 -30.220 -32.480 3549.900 ;
        RECT 121.470 -39.820 124.570 3559.500 ;
        RECT 301.470 -39.820 304.570 3559.500 ;
        RECT 481.470 760.000 484.570 3559.500 ;
        RECT 481.470 -39.820 484.570 490.000 ;
        RECT 661.470 -39.820 664.570 3559.500 ;
        RECT 841.470 -39.820 844.570 3559.500 ;
        RECT 1021.470 -39.820 1024.570 3559.500 ;
        RECT 1201.470 -39.820 1204.570 3559.500 ;
        RECT 1381.470 -39.820 1384.570 3559.500 ;
        RECT 1561.470 -39.820 1564.570 3559.500 ;
        RECT 1741.470 -39.820 1744.570 3559.500 ;
        RECT 1921.470 -39.820 1924.570 3559.500 ;
        RECT 2101.470 -39.820 2104.570 3559.500 ;
        RECT 2281.470 -39.820 2284.570 3559.500 ;
        RECT 2461.470 -39.820 2464.570 3559.500 ;
        RECT 2641.470 -39.820 2644.570 3559.500 ;
        RECT 2821.470 -39.820 2824.570 3559.500 ;
        RECT 2952.100 -30.220 2955.200 3549.900 ;
      LAYER via4 ;
        RECT -35.420 3548.560 -34.240 3549.740 ;
        RECT -33.820 3548.560 -32.640 3549.740 ;
        RECT -35.420 3546.960 -34.240 3548.140 ;
        RECT -33.820 3546.960 -32.640 3548.140 ;
        RECT -35.420 3368.590 -34.240 3369.770 ;
        RECT -33.820 3368.590 -32.640 3369.770 ;
        RECT -35.420 3366.990 -34.240 3368.170 ;
        RECT -33.820 3366.990 -32.640 3368.170 ;
        RECT -35.420 3188.590 -34.240 3189.770 ;
        RECT -33.820 3188.590 -32.640 3189.770 ;
        RECT -35.420 3186.990 -34.240 3188.170 ;
        RECT -33.820 3186.990 -32.640 3188.170 ;
        RECT -35.420 3008.590 -34.240 3009.770 ;
        RECT -33.820 3008.590 -32.640 3009.770 ;
        RECT -35.420 3006.990 -34.240 3008.170 ;
        RECT -33.820 3006.990 -32.640 3008.170 ;
        RECT -35.420 2828.590 -34.240 2829.770 ;
        RECT -33.820 2828.590 -32.640 2829.770 ;
        RECT -35.420 2826.990 -34.240 2828.170 ;
        RECT -33.820 2826.990 -32.640 2828.170 ;
        RECT -35.420 2648.590 -34.240 2649.770 ;
        RECT -33.820 2648.590 -32.640 2649.770 ;
        RECT -35.420 2646.990 -34.240 2648.170 ;
        RECT -33.820 2646.990 -32.640 2648.170 ;
        RECT -35.420 2468.590 -34.240 2469.770 ;
        RECT -33.820 2468.590 -32.640 2469.770 ;
        RECT -35.420 2466.990 -34.240 2468.170 ;
        RECT -33.820 2466.990 -32.640 2468.170 ;
        RECT -35.420 2288.590 -34.240 2289.770 ;
        RECT -33.820 2288.590 -32.640 2289.770 ;
        RECT -35.420 2286.990 -34.240 2288.170 ;
        RECT -33.820 2286.990 -32.640 2288.170 ;
        RECT -35.420 2108.590 -34.240 2109.770 ;
        RECT -33.820 2108.590 -32.640 2109.770 ;
        RECT -35.420 2106.990 -34.240 2108.170 ;
        RECT -33.820 2106.990 -32.640 2108.170 ;
        RECT -35.420 1928.590 -34.240 1929.770 ;
        RECT -33.820 1928.590 -32.640 1929.770 ;
        RECT -35.420 1926.990 -34.240 1928.170 ;
        RECT -33.820 1926.990 -32.640 1928.170 ;
        RECT -35.420 1748.590 -34.240 1749.770 ;
        RECT -33.820 1748.590 -32.640 1749.770 ;
        RECT -35.420 1746.990 -34.240 1748.170 ;
        RECT -33.820 1746.990 -32.640 1748.170 ;
        RECT -35.420 1568.590 -34.240 1569.770 ;
        RECT -33.820 1568.590 -32.640 1569.770 ;
        RECT -35.420 1566.990 -34.240 1568.170 ;
        RECT -33.820 1566.990 -32.640 1568.170 ;
        RECT -35.420 1388.590 -34.240 1389.770 ;
        RECT -33.820 1388.590 -32.640 1389.770 ;
        RECT -35.420 1386.990 -34.240 1388.170 ;
        RECT -33.820 1386.990 -32.640 1388.170 ;
        RECT -35.420 1208.590 -34.240 1209.770 ;
        RECT -33.820 1208.590 -32.640 1209.770 ;
        RECT -35.420 1206.990 -34.240 1208.170 ;
        RECT -33.820 1206.990 -32.640 1208.170 ;
        RECT -35.420 1028.590 -34.240 1029.770 ;
        RECT -33.820 1028.590 -32.640 1029.770 ;
        RECT -35.420 1026.990 -34.240 1028.170 ;
        RECT -33.820 1026.990 -32.640 1028.170 ;
        RECT -35.420 848.590 -34.240 849.770 ;
        RECT -33.820 848.590 -32.640 849.770 ;
        RECT -35.420 846.990 -34.240 848.170 ;
        RECT -33.820 846.990 -32.640 848.170 ;
        RECT -35.420 668.590 -34.240 669.770 ;
        RECT -33.820 668.590 -32.640 669.770 ;
        RECT -35.420 666.990 -34.240 668.170 ;
        RECT -33.820 666.990 -32.640 668.170 ;
        RECT -35.420 488.590 -34.240 489.770 ;
        RECT -33.820 488.590 -32.640 489.770 ;
        RECT -35.420 486.990 -34.240 488.170 ;
        RECT -33.820 486.990 -32.640 488.170 ;
        RECT -35.420 308.590 -34.240 309.770 ;
        RECT -33.820 308.590 -32.640 309.770 ;
        RECT -35.420 306.990 -34.240 308.170 ;
        RECT -33.820 306.990 -32.640 308.170 ;
        RECT -35.420 128.590 -34.240 129.770 ;
        RECT -33.820 128.590 -32.640 129.770 ;
        RECT -35.420 126.990 -34.240 128.170 ;
        RECT -33.820 126.990 -32.640 128.170 ;
        RECT -35.420 -28.460 -34.240 -27.280 ;
        RECT -33.820 -28.460 -32.640 -27.280 ;
        RECT -35.420 -30.060 -34.240 -28.880 ;
        RECT -33.820 -30.060 -32.640 -28.880 ;
        RECT 121.630 3548.560 122.810 3549.740 ;
        RECT 123.230 3548.560 124.410 3549.740 ;
        RECT 121.630 3546.960 122.810 3548.140 ;
        RECT 123.230 3546.960 124.410 3548.140 ;
        RECT 121.630 3368.590 122.810 3369.770 ;
        RECT 123.230 3368.590 124.410 3369.770 ;
        RECT 121.630 3366.990 122.810 3368.170 ;
        RECT 123.230 3366.990 124.410 3368.170 ;
        RECT 121.630 3188.590 122.810 3189.770 ;
        RECT 123.230 3188.590 124.410 3189.770 ;
        RECT 121.630 3186.990 122.810 3188.170 ;
        RECT 123.230 3186.990 124.410 3188.170 ;
        RECT 121.630 3008.590 122.810 3009.770 ;
        RECT 123.230 3008.590 124.410 3009.770 ;
        RECT 121.630 3006.990 122.810 3008.170 ;
        RECT 123.230 3006.990 124.410 3008.170 ;
        RECT 121.630 2828.590 122.810 2829.770 ;
        RECT 123.230 2828.590 124.410 2829.770 ;
        RECT 121.630 2826.990 122.810 2828.170 ;
        RECT 123.230 2826.990 124.410 2828.170 ;
        RECT 121.630 2648.590 122.810 2649.770 ;
        RECT 123.230 2648.590 124.410 2649.770 ;
        RECT 121.630 2646.990 122.810 2648.170 ;
        RECT 123.230 2646.990 124.410 2648.170 ;
        RECT 121.630 2468.590 122.810 2469.770 ;
        RECT 123.230 2468.590 124.410 2469.770 ;
        RECT 121.630 2466.990 122.810 2468.170 ;
        RECT 123.230 2466.990 124.410 2468.170 ;
        RECT 121.630 2288.590 122.810 2289.770 ;
        RECT 123.230 2288.590 124.410 2289.770 ;
        RECT 121.630 2286.990 122.810 2288.170 ;
        RECT 123.230 2286.990 124.410 2288.170 ;
        RECT 121.630 2108.590 122.810 2109.770 ;
        RECT 123.230 2108.590 124.410 2109.770 ;
        RECT 121.630 2106.990 122.810 2108.170 ;
        RECT 123.230 2106.990 124.410 2108.170 ;
        RECT 121.630 1928.590 122.810 1929.770 ;
        RECT 123.230 1928.590 124.410 1929.770 ;
        RECT 121.630 1926.990 122.810 1928.170 ;
        RECT 123.230 1926.990 124.410 1928.170 ;
        RECT 121.630 1748.590 122.810 1749.770 ;
        RECT 123.230 1748.590 124.410 1749.770 ;
        RECT 121.630 1746.990 122.810 1748.170 ;
        RECT 123.230 1746.990 124.410 1748.170 ;
        RECT 121.630 1568.590 122.810 1569.770 ;
        RECT 123.230 1568.590 124.410 1569.770 ;
        RECT 121.630 1566.990 122.810 1568.170 ;
        RECT 123.230 1566.990 124.410 1568.170 ;
        RECT 121.630 1388.590 122.810 1389.770 ;
        RECT 123.230 1388.590 124.410 1389.770 ;
        RECT 121.630 1386.990 122.810 1388.170 ;
        RECT 123.230 1386.990 124.410 1388.170 ;
        RECT 121.630 1208.590 122.810 1209.770 ;
        RECT 123.230 1208.590 124.410 1209.770 ;
        RECT 121.630 1206.990 122.810 1208.170 ;
        RECT 123.230 1206.990 124.410 1208.170 ;
        RECT 121.630 1028.590 122.810 1029.770 ;
        RECT 123.230 1028.590 124.410 1029.770 ;
        RECT 121.630 1026.990 122.810 1028.170 ;
        RECT 123.230 1026.990 124.410 1028.170 ;
        RECT 121.630 848.590 122.810 849.770 ;
        RECT 123.230 848.590 124.410 849.770 ;
        RECT 121.630 846.990 122.810 848.170 ;
        RECT 123.230 846.990 124.410 848.170 ;
        RECT 121.630 668.590 122.810 669.770 ;
        RECT 123.230 668.590 124.410 669.770 ;
        RECT 121.630 666.990 122.810 668.170 ;
        RECT 123.230 666.990 124.410 668.170 ;
        RECT 121.630 488.590 122.810 489.770 ;
        RECT 123.230 488.590 124.410 489.770 ;
        RECT 121.630 486.990 122.810 488.170 ;
        RECT 123.230 486.990 124.410 488.170 ;
        RECT 121.630 308.590 122.810 309.770 ;
        RECT 123.230 308.590 124.410 309.770 ;
        RECT 121.630 306.990 122.810 308.170 ;
        RECT 123.230 306.990 124.410 308.170 ;
        RECT 121.630 128.590 122.810 129.770 ;
        RECT 123.230 128.590 124.410 129.770 ;
        RECT 121.630 126.990 122.810 128.170 ;
        RECT 123.230 126.990 124.410 128.170 ;
        RECT 121.630 -28.460 122.810 -27.280 ;
        RECT 123.230 -28.460 124.410 -27.280 ;
        RECT 121.630 -30.060 122.810 -28.880 ;
        RECT 123.230 -30.060 124.410 -28.880 ;
        RECT 301.630 3548.560 302.810 3549.740 ;
        RECT 303.230 3548.560 304.410 3549.740 ;
        RECT 301.630 3546.960 302.810 3548.140 ;
        RECT 303.230 3546.960 304.410 3548.140 ;
        RECT 301.630 3368.590 302.810 3369.770 ;
        RECT 303.230 3368.590 304.410 3369.770 ;
        RECT 301.630 3366.990 302.810 3368.170 ;
        RECT 303.230 3366.990 304.410 3368.170 ;
        RECT 301.630 3188.590 302.810 3189.770 ;
        RECT 303.230 3188.590 304.410 3189.770 ;
        RECT 301.630 3186.990 302.810 3188.170 ;
        RECT 303.230 3186.990 304.410 3188.170 ;
        RECT 301.630 3008.590 302.810 3009.770 ;
        RECT 303.230 3008.590 304.410 3009.770 ;
        RECT 301.630 3006.990 302.810 3008.170 ;
        RECT 303.230 3006.990 304.410 3008.170 ;
        RECT 301.630 2828.590 302.810 2829.770 ;
        RECT 303.230 2828.590 304.410 2829.770 ;
        RECT 301.630 2826.990 302.810 2828.170 ;
        RECT 303.230 2826.990 304.410 2828.170 ;
        RECT 301.630 2648.590 302.810 2649.770 ;
        RECT 303.230 2648.590 304.410 2649.770 ;
        RECT 301.630 2646.990 302.810 2648.170 ;
        RECT 303.230 2646.990 304.410 2648.170 ;
        RECT 301.630 2468.590 302.810 2469.770 ;
        RECT 303.230 2468.590 304.410 2469.770 ;
        RECT 301.630 2466.990 302.810 2468.170 ;
        RECT 303.230 2466.990 304.410 2468.170 ;
        RECT 301.630 2288.590 302.810 2289.770 ;
        RECT 303.230 2288.590 304.410 2289.770 ;
        RECT 301.630 2286.990 302.810 2288.170 ;
        RECT 303.230 2286.990 304.410 2288.170 ;
        RECT 301.630 2108.590 302.810 2109.770 ;
        RECT 303.230 2108.590 304.410 2109.770 ;
        RECT 301.630 2106.990 302.810 2108.170 ;
        RECT 303.230 2106.990 304.410 2108.170 ;
        RECT 301.630 1928.590 302.810 1929.770 ;
        RECT 303.230 1928.590 304.410 1929.770 ;
        RECT 301.630 1926.990 302.810 1928.170 ;
        RECT 303.230 1926.990 304.410 1928.170 ;
        RECT 301.630 1748.590 302.810 1749.770 ;
        RECT 303.230 1748.590 304.410 1749.770 ;
        RECT 301.630 1746.990 302.810 1748.170 ;
        RECT 303.230 1746.990 304.410 1748.170 ;
        RECT 301.630 1568.590 302.810 1569.770 ;
        RECT 303.230 1568.590 304.410 1569.770 ;
        RECT 301.630 1566.990 302.810 1568.170 ;
        RECT 303.230 1566.990 304.410 1568.170 ;
        RECT 301.630 1388.590 302.810 1389.770 ;
        RECT 303.230 1388.590 304.410 1389.770 ;
        RECT 301.630 1386.990 302.810 1388.170 ;
        RECT 303.230 1386.990 304.410 1388.170 ;
        RECT 301.630 1208.590 302.810 1209.770 ;
        RECT 303.230 1208.590 304.410 1209.770 ;
        RECT 301.630 1206.990 302.810 1208.170 ;
        RECT 303.230 1206.990 304.410 1208.170 ;
        RECT 301.630 1028.590 302.810 1029.770 ;
        RECT 303.230 1028.590 304.410 1029.770 ;
        RECT 301.630 1026.990 302.810 1028.170 ;
        RECT 303.230 1026.990 304.410 1028.170 ;
        RECT 301.630 848.590 302.810 849.770 ;
        RECT 303.230 848.590 304.410 849.770 ;
        RECT 301.630 846.990 302.810 848.170 ;
        RECT 303.230 846.990 304.410 848.170 ;
        RECT 481.630 3548.560 482.810 3549.740 ;
        RECT 483.230 3548.560 484.410 3549.740 ;
        RECT 481.630 3546.960 482.810 3548.140 ;
        RECT 483.230 3546.960 484.410 3548.140 ;
        RECT 481.630 3368.590 482.810 3369.770 ;
        RECT 483.230 3368.590 484.410 3369.770 ;
        RECT 481.630 3366.990 482.810 3368.170 ;
        RECT 483.230 3366.990 484.410 3368.170 ;
        RECT 481.630 3188.590 482.810 3189.770 ;
        RECT 483.230 3188.590 484.410 3189.770 ;
        RECT 481.630 3186.990 482.810 3188.170 ;
        RECT 483.230 3186.990 484.410 3188.170 ;
        RECT 481.630 3008.590 482.810 3009.770 ;
        RECT 483.230 3008.590 484.410 3009.770 ;
        RECT 481.630 3006.990 482.810 3008.170 ;
        RECT 483.230 3006.990 484.410 3008.170 ;
        RECT 481.630 2828.590 482.810 2829.770 ;
        RECT 483.230 2828.590 484.410 2829.770 ;
        RECT 481.630 2826.990 482.810 2828.170 ;
        RECT 483.230 2826.990 484.410 2828.170 ;
        RECT 481.630 2648.590 482.810 2649.770 ;
        RECT 483.230 2648.590 484.410 2649.770 ;
        RECT 481.630 2646.990 482.810 2648.170 ;
        RECT 483.230 2646.990 484.410 2648.170 ;
        RECT 481.630 2468.590 482.810 2469.770 ;
        RECT 483.230 2468.590 484.410 2469.770 ;
        RECT 481.630 2466.990 482.810 2468.170 ;
        RECT 483.230 2466.990 484.410 2468.170 ;
        RECT 481.630 2288.590 482.810 2289.770 ;
        RECT 483.230 2288.590 484.410 2289.770 ;
        RECT 481.630 2286.990 482.810 2288.170 ;
        RECT 483.230 2286.990 484.410 2288.170 ;
        RECT 481.630 2108.590 482.810 2109.770 ;
        RECT 483.230 2108.590 484.410 2109.770 ;
        RECT 481.630 2106.990 482.810 2108.170 ;
        RECT 483.230 2106.990 484.410 2108.170 ;
        RECT 481.630 1928.590 482.810 1929.770 ;
        RECT 483.230 1928.590 484.410 1929.770 ;
        RECT 481.630 1926.990 482.810 1928.170 ;
        RECT 483.230 1926.990 484.410 1928.170 ;
        RECT 481.630 1748.590 482.810 1749.770 ;
        RECT 483.230 1748.590 484.410 1749.770 ;
        RECT 481.630 1746.990 482.810 1748.170 ;
        RECT 483.230 1746.990 484.410 1748.170 ;
        RECT 481.630 1568.590 482.810 1569.770 ;
        RECT 483.230 1568.590 484.410 1569.770 ;
        RECT 481.630 1566.990 482.810 1568.170 ;
        RECT 483.230 1566.990 484.410 1568.170 ;
        RECT 481.630 1388.590 482.810 1389.770 ;
        RECT 483.230 1388.590 484.410 1389.770 ;
        RECT 481.630 1386.990 482.810 1388.170 ;
        RECT 483.230 1386.990 484.410 1388.170 ;
        RECT 481.630 1208.590 482.810 1209.770 ;
        RECT 483.230 1208.590 484.410 1209.770 ;
        RECT 481.630 1206.990 482.810 1208.170 ;
        RECT 483.230 1206.990 484.410 1208.170 ;
        RECT 481.630 1028.590 482.810 1029.770 ;
        RECT 483.230 1028.590 484.410 1029.770 ;
        RECT 481.630 1026.990 482.810 1028.170 ;
        RECT 483.230 1026.990 484.410 1028.170 ;
        RECT 481.630 848.590 482.810 849.770 ;
        RECT 483.230 848.590 484.410 849.770 ;
        RECT 481.630 846.990 482.810 848.170 ;
        RECT 483.230 846.990 484.410 848.170 ;
        RECT 661.630 3548.560 662.810 3549.740 ;
        RECT 663.230 3548.560 664.410 3549.740 ;
        RECT 661.630 3546.960 662.810 3548.140 ;
        RECT 663.230 3546.960 664.410 3548.140 ;
        RECT 661.630 3368.590 662.810 3369.770 ;
        RECT 663.230 3368.590 664.410 3369.770 ;
        RECT 661.630 3366.990 662.810 3368.170 ;
        RECT 663.230 3366.990 664.410 3368.170 ;
        RECT 661.630 3188.590 662.810 3189.770 ;
        RECT 663.230 3188.590 664.410 3189.770 ;
        RECT 661.630 3186.990 662.810 3188.170 ;
        RECT 663.230 3186.990 664.410 3188.170 ;
        RECT 661.630 3008.590 662.810 3009.770 ;
        RECT 663.230 3008.590 664.410 3009.770 ;
        RECT 661.630 3006.990 662.810 3008.170 ;
        RECT 663.230 3006.990 664.410 3008.170 ;
        RECT 661.630 2828.590 662.810 2829.770 ;
        RECT 663.230 2828.590 664.410 2829.770 ;
        RECT 661.630 2826.990 662.810 2828.170 ;
        RECT 663.230 2826.990 664.410 2828.170 ;
        RECT 661.630 2648.590 662.810 2649.770 ;
        RECT 663.230 2648.590 664.410 2649.770 ;
        RECT 661.630 2646.990 662.810 2648.170 ;
        RECT 663.230 2646.990 664.410 2648.170 ;
        RECT 661.630 2468.590 662.810 2469.770 ;
        RECT 663.230 2468.590 664.410 2469.770 ;
        RECT 661.630 2466.990 662.810 2468.170 ;
        RECT 663.230 2466.990 664.410 2468.170 ;
        RECT 661.630 2288.590 662.810 2289.770 ;
        RECT 663.230 2288.590 664.410 2289.770 ;
        RECT 661.630 2286.990 662.810 2288.170 ;
        RECT 663.230 2286.990 664.410 2288.170 ;
        RECT 661.630 2108.590 662.810 2109.770 ;
        RECT 663.230 2108.590 664.410 2109.770 ;
        RECT 661.630 2106.990 662.810 2108.170 ;
        RECT 663.230 2106.990 664.410 2108.170 ;
        RECT 661.630 1928.590 662.810 1929.770 ;
        RECT 663.230 1928.590 664.410 1929.770 ;
        RECT 661.630 1926.990 662.810 1928.170 ;
        RECT 663.230 1926.990 664.410 1928.170 ;
        RECT 661.630 1748.590 662.810 1749.770 ;
        RECT 663.230 1748.590 664.410 1749.770 ;
        RECT 661.630 1746.990 662.810 1748.170 ;
        RECT 663.230 1746.990 664.410 1748.170 ;
        RECT 661.630 1568.590 662.810 1569.770 ;
        RECT 663.230 1568.590 664.410 1569.770 ;
        RECT 661.630 1566.990 662.810 1568.170 ;
        RECT 663.230 1566.990 664.410 1568.170 ;
        RECT 661.630 1388.590 662.810 1389.770 ;
        RECT 663.230 1388.590 664.410 1389.770 ;
        RECT 661.630 1386.990 662.810 1388.170 ;
        RECT 663.230 1386.990 664.410 1388.170 ;
        RECT 661.630 1208.590 662.810 1209.770 ;
        RECT 663.230 1208.590 664.410 1209.770 ;
        RECT 661.630 1206.990 662.810 1208.170 ;
        RECT 663.230 1206.990 664.410 1208.170 ;
        RECT 661.630 1028.590 662.810 1029.770 ;
        RECT 663.230 1028.590 664.410 1029.770 ;
        RECT 661.630 1026.990 662.810 1028.170 ;
        RECT 663.230 1026.990 664.410 1028.170 ;
        RECT 661.630 848.590 662.810 849.770 ;
        RECT 663.230 848.590 664.410 849.770 ;
        RECT 661.630 846.990 662.810 848.170 ;
        RECT 663.230 846.990 664.410 848.170 ;
        RECT 301.630 668.590 302.810 669.770 ;
        RECT 303.230 668.590 304.410 669.770 ;
        RECT 301.630 666.990 302.810 668.170 ;
        RECT 303.230 666.990 304.410 668.170 ;
        RECT 661.630 668.590 662.810 669.770 ;
        RECT 663.230 668.590 664.410 669.770 ;
        RECT 661.630 666.990 662.810 668.170 ;
        RECT 663.230 666.990 664.410 668.170 ;
        RECT 301.630 488.590 302.810 489.770 ;
        RECT 303.230 488.590 304.410 489.770 ;
        RECT 301.630 486.990 302.810 488.170 ;
        RECT 303.230 486.990 304.410 488.170 ;
        RECT 301.630 308.590 302.810 309.770 ;
        RECT 303.230 308.590 304.410 309.770 ;
        RECT 301.630 306.990 302.810 308.170 ;
        RECT 303.230 306.990 304.410 308.170 ;
        RECT 301.630 128.590 302.810 129.770 ;
        RECT 303.230 128.590 304.410 129.770 ;
        RECT 301.630 126.990 302.810 128.170 ;
        RECT 303.230 126.990 304.410 128.170 ;
        RECT 301.630 -28.460 302.810 -27.280 ;
        RECT 303.230 -28.460 304.410 -27.280 ;
        RECT 301.630 -30.060 302.810 -28.880 ;
        RECT 303.230 -30.060 304.410 -28.880 ;
        RECT 481.630 488.590 482.810 489.770 ;
        RECT 483.230 488.590 484.410 489.770 ;
        RECT 481.630 486.990 482.810 488.170 ;
        RECT 483.230 486.990 484.410 488.170 ;
        RECT 481.630 308.590 482.810 309.770 ;
        RECT 483.230 308.590 484.410 309.770 ;
        RECT 481.630 306.990 482.810 308.170 ;
        RECT 483.230 306.990 484.410 308.170 ;
        RECT 481.630 128.590 482.810 129.770 ;
        RECT 483.230 128.590 484.410 129.770 ;
        RECT 481.630 126.990 482.810 128.170 ;
        RECT 483.230 126.990 484.410 128.170 ;
        RECT 481.630 -28.460 482.810 -27.280 ;
        RECT 483.230 -28.460 484.410 -27.280 ;
        RECT 481.630 -30.060 482.810 -28.880 ;
        RECT 483.230 -30.060 484.410 -28.880 ;
        RECT 661.630 488.590 662.810 489.770 ;
        RECT 663.230 488.590 664.410 489.770 ;
        RECT 661.630 486.990 662.810 488.170 ;
        RECT 663.230 486.990 664.410 488.170 ;
        RECT 661.630 308.590 662.810 309.770 ;
        RECT 663.230 308.590 664.410 309.770 ;
        RECT 661.630 306.990 662.810 308.170 ;
        RECT 663.230 306.990 664.410 308.170 ;
        RECT 661.630 128.590 662.810 129.770 ;
        RECT 663.230 128.590 664.410 129.770 ;
        RECT 661.630 126.990 662.810 128.170 ;
        RECT 663.230 126.990 664.410 128.170 ;
        RECT 661.630 -28.460 662.810 -27.280 ;
        RECT 663.230 -28.460 664.410 -27.280 ;
        RECT 661.630 -30.060 662.810 -28.880 ;
        RECT 663.230 -30.060 664.410 -28.880 ;
        RECT 841.630 3548.560 842.810 3549.740 ;
        RECT 843.230 3548.560 844.410 3549.740 ;
        RECT 841.630 3546.960 842.810 3548.140 ;
        RECT 843.230 3546.960 844.410 3548.140 ;
        RECT 841.630 3368.590 842.810 3369.770 ;
        RECT 843.230 3368.590 844.410 3369.770 ;
        RECT 841.630 3366.990 842.810 3368.170 ;
        RECT 843.230 3366.990 844.410 3368.170 ;
        RECT 841.630 3188.590 842.810 3189.770 ;
        RECT 843.230 3188.590 844.410 3189.770 ;
        RECT 841.630 3186.990 842.810 3188.170 ;
        RECT 843.230 3186.990 844.410 3188.170 ;
        RECT 841.630 3008.590 842.810 3009.770 ;
        RECT 843.230 3008.590 844.410 3009.770 ;
        RECT 841.630 3006.990 842.810 3008.170 ;
        RECT 843.230 3006.990 844.410 3008.170 ;
        RECT 841.630 2828.590 842.810 2829.770 ;
        RECT 843.230 2828.590 844.410 2829.770 ;
        RECT 841.630 2826.990 842.810 2828.170 ;
        RECT 843.230 2826.990 844.410 2828.170 ;
        RECT 841.630 2648.590 842.810 2649.770 ;
        RECT 843.230 2648.590 844.410 2649.770 ;
        RECT 841.630 2646.990 842.810 2648.170 ;
        RECT 843.230 2646.990 844.410 2648.170 ;
        RECT 841.630 2468.590 842.810 2469.770 ;
        RECT 843.230 2468.590 844.410 2469.770 ;
        RECT 841.630 2466.990 842.810 2468.170 ;
        RECT 843.230 2466.990 844.410 2468.170 ;
        RECT 841.630 2288.590 842.810 2289.770 ;
        RECT 843.230 2288.590 844.410 2289.770 ;
        RECT 841.630 2286.990 842.810 2288.170 ;
        RECT 843.230 2286.990 844.410 2288.170 ;
        RECT 841.630 2108.590 842.810 2109.770 ;
        RECT 843.230 2108.590 844.410 2109.770 ;
        RECT 841.630 2106.990 842.810 2108.170 ;
        RECT 843.230 2106.990 844.410 2108.170 ;
        RECT 841.630 1928.590 842.810 1929.770 ;
        RECT 843.230 1928.590 844.410 1929.770 ;
        RECT 841.630 1926.990 842.810 1928.170 ;
        RECT 843.230 1926.990 844.410 1928.170 ;
        RECT 841.630 1748.590 842.810 1749.770 ;
        RECT 843.230 1748.590 844.410 1749.770 ;
        RECT 841.630 1746.990 842.810 1748.170 ;
        RECT 843.230 1746.990 844.410 1748.170 ;
        RECT 841.630 1568.590 842.810 1569.770 ;
        RECT 843.230 1568.590 844.410 1569.770 ;
        RECT 841.630 1566.990 842.810 1568.170 ;
        RECT 843.230 1566.990 844.410 1568.170 ;
        RECT 841.630 1388.590 842.810 1389.770 ;
        RECT 843.230 1388.590 844.410 1389.770 ;
        RECT 841.630 1386.990 842.810 1388.170 ;
        RECT 843.230 1386.990 844.410 1388.170 ;
        RECT 841.630 1208.590 842.810 1209.770 ;
        RECT 843.230 1208.590 844.410 1209.770 ;
        RECT 841.630 1206.990 842.810 1208.170 ;
        RECT 843.230 1206.990 844.410 1208.170 ;
        RECT 841.630 1028.590 842.810 1029.770 ;
        RECT 843.230 1028.590 844.410 1029.770 ;
        RECT 841.630 1026.990 842.810 1028.170 ;
        RECT 843.230 1026.990 844.410 1028.170 ;
        RECT 841.630 848.590 842.810 849.770 ;
        RECT 843.230 848.590 844.410 849.770 ;
        RECT 841.630 846.990 842.810 848.170 ;
        RECT 843.230 846.990 844.410 848.170 ;
        RECT 841.630 668.590 842.810 669.770 ;
        RECT 843.230 668.590 844.410 669.770 ;
        RECT 841.630 666.990 842.810 668.170 ;
        RECT 843.230 666.990 844.410 668.170 ;
        RECT 841.630 488.590 842.810 489.770 ;
        RECT 843.230 488.590 844.410 489.770 ;
        RECT 841.630 486.990 842.810 488.170 ;
        RECT 843.230 486.990 844.410 488.170 ;
        RECT 841.630 308.590 842.810 309.770 ;
        RECT 843.230 308.590 844.410 309.770 ;
        RECT 841.630 306.990 842.810 308.170 ;
        RECT 843.230 306.990 844.410 308.170 ;
        RECT 841.630 128.590 842.810 129.770 ;
        RECT 843.230 128.590 844.410 129.770 ;
        RECT 841.630 126.990 842.810 128.170 ;
        RECT 843.230 126.990 844.410 128.170 ;
        RECT 841.630 -28.460 842.810 -27.280 ;
        RECT 843.230 -28.460 844.410 -27.280 ;
        RECT 841.630 -30.060 842.810 -28.880 ;
        RECT 843.230 -30.060 844.410 -28.880 ;
        RECT 1021.630 3548.560 1022.810 3549.740 ;
        RECT 1023.230 3548.560 1024.410 3549.740 ;
        RECT 1021.630 3546.960 1022.810 3548.140 ;
        RECT 1023.230 3546.960 1024.410 3548.140 ;
        RECT 1021.630 3368.590 1022.810 3369.770 ;
        RECT 1023.230 3368.590 1024.410 3369.770 ;
        RECT 1021.630 3366.990 1022.810 3368.170 ;
        RECT 1023.230 3366.990 1024.410 3368.170 ;
        RECT 1021.630 3188.590 1022.810 3189.770 ;
        RECT 1023.230 3188.590 1024.410 3189.770 ;
        RECT 1021.630 3186.990 1022.810 3188.170 ;
        RECT 1023.230 3186.990 1024.410 3188.170 ;
        RECT 1021.630 3008.590 1022.810 3009.770 ;
        RECT 1023.230 3008.590 1024.410 3009.770 ;
        RECT 1021.630 3006.990 1022.810 3008.170 ;
        RECT 1023.230 3006.990 1024.410 3008.170 ;
        RECT 1021.630 2828.590 1022.810 2829.770 ;
        RECT 1023.230 2828.590 1024.410 2829.770 ;
        RECT 1021.630 2826.990 1022.810 2828.170 ;
        RECT 1023.230 2826.990 1024.410 2828.170 ;
        RECT 1021.630 2648.590 1022.810 2649.770 ;
        RECT 1023.230 2648.590 1024.410 2649.770 ;
        RECT 1021.630 2646.990 1022.810 2648.170 ;
        RECT 1023.230 2646.990 1024.410 2648.170 ;
        RECT 1021.630 2468.590 1022.810 2469.770 ;
        RECT 1023.230 2468.590 1024.410 2469.770 ;
        RECT 1021.630 2466.990 1022.810 2468.170 ;
        RECT 1023.230 2466.990 1024.410 2468.170 ;
        RECT 1021.630 2288.590 1022.810 2289.770 ;
        RECT 1023.230 2288.590 1024.410 2289.770 ;
        RECT 1021.630 2286.990 1022.810 2288.170 ;
        RECT 1023.230 2286.990 1024.410 2288.170 ;
        RECT 1021.630 2108.590 1022.810 2109.770 ;
        RECT 1023.230 2108.590 1024.410 2109.770 ;
        RECT 1021.630 2106.990 1022.810 2108.170 ;
        RECT 1023.230 2106.990 1024.410 2108.170 ;
        RECT 1021.630 1928.590 1022.810 1929.770 ;
        RECT 1023.230 1928.590 1024.410 1929.770 ;
        RECT 1021.630 1926.990 1022.810 1928.170 ;
        RECT 1023.230 1926.990 1024.410 1928.170 ;
        RECT 1021.630 1748.590 1022.810 1749.770 ;
        RECT 1023.230 1748.590 1024.410 1749.770 ;
        RECT 1021.630 1746.990 1022.810 1748.170 ;
        RECT 1023.230 1746.990 1024.410 1748.170 ;
        RECT 1021.630 1568.590 1022.810 1569.770 ;
        RECT 1023.230 1568.590 1024.410 1569.770 ;
        RECT 1021.630 1566.990 1022.810 1568.170 ;
        RECT 1023.230 1566.990 1024.410 1568.170 ;
        RECT 1021.630 1388.590 1022.810 1389.770 ;
        RECT 1023.230 1388.590 1024.410 1389.770 ;
        RECT 1021.630 1386.990 1022.810 1388.170 ;
        RECT 1023.230 1386.990 1024.410 1388.170 ;
        RECT 1021.630 1208.590 1022.810 1209.770 ;
        RECT 1023.230 1208.590 1024.410 1209.770 ;
        RECT 1021.630 1206.990 1022.810 1208.170 ;
        RECT 1023.230 1206.990 1024.410 1208.170 ;
        RECT 1021.630 1028.590 1022.810 1029.770 ;
        RECT 1023.230 1028.590 1024.410 1029.770 ;
        RECT 1021.630 1026.990 1022.810 1028.170 ;
        RECT 1023.230 1026.990 1024.410 1028.170 ;
        RECT 1021.630 848.590 1022.810 849.770 ;
        RECT 1023.230 848.590 1024.410 849.770 ;
        RECT 1021.630 846.990 1022.810 848.170 ;
        RECT 1023.230 846.990 1024.410 848.170 ;
        RECT 1021.630 668.590 1022.810 669.770 ;
        RECT 1023.230 668.590 1024.410 669.770 ;
        RECT 1021.630 666.990 1022.810 668.170 ;
        RECT 1023.230 666.990 1024.410 668.170 ;
        RECT 1021.630 488.590 1022.810 489.770 ;
        RECT 1023.230 488.590 1024.410 489.770 ;
        RECT 1021.630 486.990 1022.810 488.170 ;
        RECT 1023.230 486.990 1024.410 488.170 ;
        RECT 1021.630 308.590 1022.810 309.770 ;
        RECT 1023.230 308.590 1024.410 309.770 ;
        RECT 1021.630 306.990 1022.810 308.170 ;
        RECT 1023.230 306.990 1024.410 308.170 ;
        RECT 1021.630 128.590 1022.810 129.770 ;
        RECT 1023.230 128.590 1024.410 129.770 ;
        RECT 1021.630 126.990 1022.810 128.170 ;
        RECT 1023.230 126.990 1024.410 128.170 ;
        RECT 1021.630 -28.460 1022.810 -27.280 ;
        RECT 1023.230 -28.460 1024.410 -27.280 ;
        RECT 1021.630 -30.060 1022.810 -28.880 ;
        RECT 1023.230 -30.060 1024.410 -28.880 ;
        RECT 1201.630 3548.560 1202.810 3549.740 ;
        RECT 1203.230 3548.560 1204.410 3549.740 ;
        RECT 1201.630 3546.960 1202.810 3548.140 ;
        RECT 1203.230 3546.960 1204.410 3548.140 ;
        RECT 1201.630 3368.590 1202.810 3369.770 ;
        RECT 1203.230 3368.590 1204.410 3369.770 ;
        RECT 1201.630 3366.990 1202.810 3368.170 ;
        RECT 1203.230 3366.990 1204.410 3368.170 ;
        RECT 1201.630 3188.590 1202.810 3189.770 ;
        RECT 1203.230 3188.590 1204.410 3189.770 ;
        RECT 1201.630 3186.990 1202.810 3188.170 ;
        RECT 1203.230 3186.990 1204.410 3188.170 ;
        RECT 1201.630 3008.590 1202.810 3009.770 ;
        RECT 1203.230 3008.590 1204.410 3009.770 ;
        RECT 1201.630 3006.990 1202.810 3008.170 ;
        RECT 1203.230 3006.990 1204.410 3008.170 ;
        RECT 1201.630 2828.590 1202.810 2829.770 ;
        RECT 1203.230 2828.590 1204.410 2829.770 ;
        RECT 1201.630 2826.990 1202.810 2828.170 ;
        RECT 1203.230 2826.990 1204.410 2828.170 ;
        RECT 1201.630 2648.590 1202.810 2649.770 ;
        RECT 1203.230 2648.590 1204.410 2649.770 ;
        RECT 1201.630 2646.990 1202.810 2648.170 ;
        RECT 1203.230 2646.990 1204.410 2648.170 ;
        RECT 1201.630 2468.590 1202.810 2469.770 ;
        RECT 1203.230 2468.590 1204.410 2469.770 ;
        RECT 1201.630 2466.990 1202.810 2468.170 ;
        RECT 1203.230 2466.990 1204.410 2468.170 ;
        RECT 1201.630 2288.590 1202.810 2289.770 ;
        RECT 1203.230 2288.590 1204.410 2289.770 ;
        RECT 1201.630 2286.990 1202.810 2288.170 ;
        RECT 1203.230 2286.990 1204.410 2288.170 ;
        RECT 1201.630 2108.590 1202.810 2109.770 ;
        RECT 1203.230 2108.590 1204.410 2109.770 ;
        RECT 1201.630 2106.990 1202.810 2108.170 ;
        RECT 1203.230 2106.990 1204.410 2108.170 ;
        RECT 1201.630 1928.590 1202.810 1929.770 ;
        RECT 1203.230 1928.590 1204.410 1929.770 ;
        RECT 1201.630 1926.990 1202.810 1928.170 ;
        RECT 1203.230 1926.990 1204.410 1928.170 ;
        RECT 1201.630 1748.590 1202.810 1749.770 ;
        RECT 1203.230 1748.590 1204.410 1749.770 ;
        RECT 1201.630 1746.990 1202.810 1748.170 ;
        RECT 1203.230 1746.990 1204.410 1748.170 ;
        RECT 1201.630 1568.590 1202.810 1569.770 ;
        RECT 1203.230 1568.590 1204.410 1569.770 ;
        RECT 1201.630 1566.990 1202.810 1568.170 ;
        RECT 1203.230 1566.990 1204.410 1568.170 ;
        RECT 1201.630 1388.590 1202.810 1389.770 ;
        RECT 1203.230 1388.590 1204.410 1389.770 ;
        RECT 1201.630 1386.990 1202.810 1388.170 ;
        RECT 1203.230 1386.990 1204.410 1388.170 ;
        RECT 1201.630 1208.590 1202.810 1209.770 ;
        RECT 1203.230 1208.590 1204.410 1209.770 ;
        RECT 1201.630 1206.990 1202.810 1208.170 ;
        RECT 1203.230 1206.990 1204.410 1208.170 ;
        RECT 1201.630 1028.590 1202.810 1029.770 ;
        RECT 1203.230 1028.590 1204.410 1029.770 ;
        RECT 1201.630 1026.990 1202.810 1028.170 ;
        RECT 1203.230 1026.990 1204.410 1028.170 ;
        RECT 1201.630 848.590 1202.810 849.770 ;
        RECT 1203.230 848.590 1204.410 849.770 ;
        RECT 1201.630 846.990 1202.810 848.170 ;
        RECT 1203.230 846.990 1204.410 848.170 ;
        RECT 1201.630 668.590 1202.810 669.770 ;
        RECT 1203.230 668.590 1204.410 669.770 ;
        RECT 1201.630 666.990 1202.810 668.170 ;
        RECT 1203.230 666.990 1204.410 668.170 ;
        RECT 1201.630 488.590 1202.810 489.770 ;
        RECT 1203.230 488.590 1204.410 489.770 ;
        RECT 1201.630 486.990 1202.810 488.170 ;
        RECT 1203.230 486.990 1204.410 488.170 ;
        RECT 1201.630 308.590 1202.810 309.770 ;
        RECT 1203.230 308.590 1204.410 309.770 ;
        RECT 1201.630 306.990 1202.810 308.170 ;
        RECT 1203.230 306.990 1204.410 308.170 ;
        RECT 1201.630 128.590 1202.810 129.770 ;
        RECT 1203.230 128.590 1204.410 129.770 ;
        RECT 1201.630 126.990 1202.810 128.170 ;
        RECT 1203.230 126.990 1204.410 128.170 ;
        RECT 1201.630 -28.460 1202.810 -27.280 ;
        RECT 1203.230 -28.460 1204.410 -27.280 ;
        RECT 1201.630 -30.060 1202.810 -28.880 ;
        RECT 1203.230 -30.060 1204.410 -28.880 ;
        RECT 1381.630 3548.560 1382.810 3549.740 ;
        RECT 1383.230 3548.560 1384.410 3549.740 ;
        RECT 1381.630 3546.960 1382.810 3548.140 ;
        RECT 1383.230 3546.960 1384.410 3548.140 ;
        RECT 1381.630 3368.590 1382.810 3369.770 ;
        RECT 1383.230 3368.590 1384.410 3369.770 ;
        RECT 1381.630 3366.990 1382.810 3368.170 ;
        RECT 1383.230 3366.990 1384.410 3368.170 ;
        RECT 1381.630 3188.590 1382.810 3189.770 ;
        RECT 1383.230 3188.590 1384.410 3189.770 ;
        RECT 1381.630 3186.990 1382.810 3188.170 ;
        RECT 1383.230 3186.990 1384.410 3188.170 ;
        RECT 1381.630 3008.590 1382.810 3009.770 ;
        RECT 1383.230 3008.590 1384.410 3009.770 ;
        RECT 1381.630 3006.990 1382.810 3008.170 ;
        RECT 1383.230 3006.990 1384.410 3008.170 ;
        RECT 1381.630 2828.590 1382.810 2829.770 ;
        RECT 1383.230 2828.590 1384.410 2829.770 ;
        RECT 1381.630 2826.990 1382.810 2828.170 ;
        RECT 1383.230 2826.990 1384.410 2828.170 ;
        RECT 1381.630 2648.590 1382.810 2649.770 ;
        RECT 1383.230 2648.590 1384.410 2649.770 ;
        RECT 1381.630 2646.990 1382.810 2648.170 ;
        RECT 1383.230 2646.990 1384.410 2648.170 ;
        RECT 1381.630 2468.590 1382.810 2469.770 ;
        RECT 1383.230 2468.590 1384.410 2469.770 ;
        RECT 1381.630 2466.990 1382.810 2468.170 ;
        RECT 1383.230 2466.990 1384.410 2468.170 ;
        RECT 1381.630 2288.590 1382.810 2289.770 ;
        RECT 1383.230 2288.590 1384.410 2289.770 ;
        RECT 1381.630 2286.990 1382.810 2288.170 ;
        RECT 1383.230 2286.990 1384.410 2288.170 ;
        RECT 1381.630 2108.590 1382.810 2109.770 ;
        RECT 1383.230 2108.590 1384.410 2109.770 ;
        RECT 1381.630 2106.990 1382.810 2108.170 ;
        RECT 1383.230 2106.990 1384.410 2108.170 ;
        RECT 1381.630 1928.590 1382.810 1929.770 ;
        RECT 1383.230 1928.590 1384.410 1929.770 ;
        RECT 1381.630 1926.990 1382.810 1928.170 ;
        RECT 1383.230 1926.990 1384.410 1928.170 ;
        RECT 1381.630 1748.590 1382.810 1749.770 ;
        RECT 1383.230 1748.590 1384.410 1749.770 ;
        RECT 1381.630 1746.990 1382.810 1748.170 ;
        RECT 1383.230 1746.990 1384.410 1748.170 ;
        RECT 1381.630 1568.590 1382.810 1569.770 ;
        RECT 1383.230 1568.590 1384.410 1569.770 ;
        RECT 1381.630 1566.990 1382.810 1568.170 ;
        RECT 1383.230 1566.990 1384.410 1568.170 ;
        RECT 1381.630 1388.590 1382.810 1389.770 ;
        RECT 1383.230 1388.590 1384.410 1389.770 ;
        RECT 1381.630 1386.990 1382.810 1388.170 ;
        RECT 1383.230 1386.990 1384.410 1388.170 ;
        RECT 1381.630 1208.590 1382.810 1209.770 ;
        RECT 1383.230 1208.590 1384.410 1209.770 ;
        RECT 1381.630 1206.990 1382.810 1208.170 ;
        RECT 1383.230 1206.990 1384.410 1208.170 ;
        RECT 1381.630 1028.590 1382.810 1029.770 ;
        RECT 1383.230 1028.590 1384.410 1029.770 ;
        RECT 1381.630 1026.990 1382.810 1028.170 ;
        RECT 1383.230 1026.990 1384.410 1028.170 ;
        RECT 1381.630 848.590 1382.810 849.770 ;
        RECT 1383.230 848.590 1384.410 849.770 ;
        RECT 1381.630 846.990 1382.810 848.170 ;
        RECT 1383.230 846.990 1384.410 848.170 ;
        RECT 1381.630 668.590 1382.810 669.770 ;
        RECT 1383.230 668.590 1384.410 669.770 ;
        RECT 1381.630 666.990 1382.810 668.170 ;
        RECT 1383.230 666.990 1384.410 668.170 ;
        RECT 1381.630 488.590 1382.810 489.770 ;
        RECT 1383.230 488.590 1384.410 489.770 ;
        RECT 1381.630 486.990 1382.810 488.170 ;
        RECT 1383.230 486.990 1384.410 488.170 ;
        RECT 1381.630 308.590 1382.810 309.770 ;
        RECT 1383.230 308.590 1384.410 309.770 ;
        RECT 1381.630 306.990 1382.810 308.170 ;
        RECT 1383.230 306.990 1384.410 308.170 ;
        RECT 1381.630 128.590 1382.810 129.770 ;
        RECT 1383.230 128.590 1384.410 129.770 ;
        RECT 1381.630 126.990 1382.810 128.170 ;
        RECT 1383.230 126.990 1384.410 128.170 ;
        RECT 1381.630 -28.460 1382.810 -27.280 ;
        RECT 1383.230 -28.460 1384.410 -27.280 ;
        RECT 1381.630 -30.060 1382.810 -28.880 ;
        RECT 1383.230 -30.060 1384.410 -28.880 ;
        RECT 1561.630 3548.560 1562.810 3549.740 ;
        RECT 1563.230 3548.560 1564.410 3549.740 ;
        RECT 1561.630 3546.960 1562.810 3548.140 ;
        RECT 1563.230 3546.960 1564.410 3548.140 ;
        RECT 1561.630 3368.590 1562.810 3369.770 ;
        RECT 1563.230 3368.590 1564.410 3369.770 ;
        RECT 1561.630 3366.990 1562.810 3368.170 ;
        RECT 1563.230 3366.990 1564.410 3368.170 ;
        RECT 1561.630 3188.590 1562.810 3189.770 ;
        RECT 1563.230 3188.590 1564.410 3189.770 ;
        RECT 1561.630 3186.990 1562.810 3188.170 ;
        RECT 1563.230 3186.990 1564.410 3188.170 ;
        RECT 1561.630 3008.590 1562.810 3009.770 ;
        RECT 1563.230 3008.590 1564.410 3009.770 ;
        RECT 1561.630 3006.990 1562.810 3008.170 ;
        RECT 1563.230 3006.990 1564.410 3008.170 ;
        RECT 1561.630 2828.590 1562.810 2829.770 ;
        RECT 1563.230 2828.590 1564.410 2829.770 ;
        RECT 1561.630 2826.990 1562.810 2828.170 ;
        RECT 1563.230 2826.990 1564.410 2828.170 ;
        RECT 1561.630 2648.590 1562.810 2649.770 ;
        RECT 1563.230 2648.590 1564.410 2649.770 ;
        RECT 1561.630 2646.990 1562.810 2648.170 ;
        RECT 1563.230 2646.990 1564.410 2648.170 ;
        RECT 1561.630 2468.590 1562.810 2469.770 ;
        RECT 1563.230 2468.590 1564.410 2469.770 ;
        RECT 1561.630 2466.990 1562.810 2468.170 ;
        RECT 1563.230 2466.990 1564.410 2468.170 ;
        RECT 1561.630 2288.590 1562.810 2289.770 ;
        RECT 1563.230 2288.590 1564.410 2289.770 ;
        RECT 1561.630 2286.990 1562.810 2288.170 ;
        RECT 1563.230 2286.990 1564.410 2288.170 ;
        RECT 1561.630 2108.590 1562.810 2109.770 ;
        RECT 1563.230 2108.590 1564.410 2109.770 ;
        RECT 1561.630 2106.990 1562.810 2108.170 ;
        RECT 1563.230 2106.990 1564.410 2108.170 ;
        RECT 1561.630 1928.590 1562.810 1929.770 ;
        RECT 1563.230 1928.590 1564.410 1929.770 ;
        RECT 1561.630 1926.990 1562.810 1928.170 ;
        RECT 1563.230 1926.990 1564.410 1928.170 ;
        RECT 1561.630 1748.590 1562.810 1749.770 ;
        RECT 1563.230 1748.590 1564.410 1749.770 ;
        RECT 1561.630 1746.990 1562.810 1748.170 ;
        RECT 1563.230 1746.990 1564.410 1748.170 ;
        RECT 1561.630 1568.590 1562.810 1569.770 ;
        RECT 1563.230 1568.590 1564.410 1569.770 ;
        RECT 1561.630 1566.990 1562.810 1568.170 ;
        RECT 1563.230 1566.990 1564.410 1568.170 ;
        RECT 1561.630 1388.590 1562.810 1389.770 ;
        RECT 1563.230 1388.590 1564.410 1389.770 ;
        RECT 1561.630 1386.990 1562.810 1388.170 ;
        RECT 1563.230 1386.990 1564.410 1388.170 ;
        RECT 1561.630 1208.590 1562.810 1209.770 ;
        RECT 1563.230 1208.590 1564.410 1209.770 ;
        RECT 1561.630 1206.990 1562.810 1208.170 ;
        RECT 1563.230 1206.990 1564.410 1208.170 ;
        RECT 1561.630 1028.590 1562.810 1029.770 ;
        RECT 1563.230 1028.590 1564.410 1029.770 ;
        RECT 1561.630 1026.990 1562.810 1028.170 ;
        RECT 1563.230 1026.990 1564.410 1028.170 ;
        RECT 1561.630 848.590 1562.810 849.770 ;
        RECT 1563.230 848.590 1564.410 849.770 ;
        RECT 1561.630 846.990 1562.810 848.170 ;
        RECT 1563.230 846.990 1564.410 848.170 ;
        RECT 1561.630 668.590 1562.810 669.770 ;
        RECT 1563.230 668.590 1564.410 669.770 ;
        RECT 1561.630 666.990 1562.810 668.170 ;
        RECT 1563.230 666.990 1564.410 668.170 ;
        RECT 1561.630 488.590 1562.810 489.770 ;
        RECT 1563.230 488.590 1564.410 489.770 ;
        RECT 1561.630 486.990 1562.810 488.170 ;
        RECT 1563.230 486.990 1564.410 488.170 ;
        RECT 1561.630 308.590 1562.810 309.770 ;
        RECT 1563.230 308.590 1564.410 309.770 ;
        RECT 1561.630 306.990 1562.810 308.170 ;
        RECT 1563.230 306.990 1564.410 308.170 ;
        RECT 1561.630 128.590 1562.810 129.770 ;
        RECT 1563.230 128.590 1564.410 129.770 ;
        RECT 1561.630 126.990 1562.810 128.170 ;
        RECT 1563.230 126.990 1564.410 128.170 ;
        RECT 1561.630 -28.460 1562.810 -27.280 ;
        RECT 1563.230 -28.460 1564.410 -27.280 ;
        RECT 1561.630 -30.060 1562.810 -28.880 ;
        RECT 1563.230 -30.060 1564.410 -28.880 ;
        RECT 1741.630 3548.560 1742.810 3549.740 ;
        RECT 1743.230 3548.560 1744.410 3549.740 ;
        RECT 1741.630 3546.960 1742.810 3548.140 ;
        RECT 1743.230 3546.960 1744.410 3548.140 ;
        RECT 1741.630 3368.590 1742.810 3369.770 ;
        RECT 1743.230 3368.590 1744.410 3369.770 ;
        RECT 1741.630 3366.990 1742.810 3368.170 ;
        RECT 1743.230 3366.990 1744.410 3368.170 ;
        RECT 1741.630 3188.590 1742.810 3189.770 ;
        RECT 1743.230 3188.590 1744.410 3189.770 ;
        RECT 1741.630 3186.990 1742.810 3188.170 ;
        RECT 1743.230 3186.990 1744.410 3188.170 ;
        RECT 1741.630 3008.590 1742.810 3009.770 ;
        RECT 1743.230 3008.590 1744.410 3009.770 ;
        RECT 1741.630 3006.990 1742.810 3008.170 ;
        RECT 1743.230 3006.990 1744.410 3008.170 ;
        RECT 1741.630 2828.590 1742.810 2829.770 ;
        RECT 1743.230 2828.590 1744.410 2829.770 ;
        RECT 1741.630 2826.990 1742.810 2828.170 ;
        RECT 1743.230 2826.990 1744.410 2828.170 ;
        RECT 1741.630 2648.590 1742.810 2649.770 ;
        RECT 1743.230 2648.590 1744.410 2649.770 ;
        RECT 1741.630 2646.990 1742.810 2648.170 ;
        RECT 1743.230 2646.990 1744.410 2648.170 ;
        RECT 1741.630 2468.590 1742.810 2469.770 ;
        RECT 1743.230 2468.590 1744.410 2469.770 ;
        RECT 1741.630 2466.990 1742.810 2468.170 ;
        RECT 1743.230 2466.990 1744.410 2468.170 ;
        RECT 1741.630 2288.590 1742.810 2289.770 ;
        RECT 1743.230 2288.590 1744.410 2289.770 ;
        RECT 1741.630 2286.990 1742.810 2288.170 ;
        RECT 1743.230 2286.990 1744.410 2288.170 ;
        RECT 1741.630 2108.590 1742.810 2109.770 ;
        RECT 1743.230 2108.590 1744.410 2109.770 ;
        RECT 1741.630 2106.990 1742.810 2108.170 ;
        RECT 1743.230 2106.990 1744.410 2108.170 ;
        RECT 1741.630 1928.590 1742.810 1929.770 ;
        RECT 1743.230 1928.590 1744.410 1929.770 ;
        RECT 1741.630 1926.990 1742.810 1928.170 ;
        RECT 1743.230 1926.990 1744.410 1928.170 ;
        RECT 1741.630 1748.590 1742.810 1749.770 ;
        RECT 1743.230 1748.590 1744.410 1749.770 ;
        RECT 1741.630 1746.990 1742.810 1748.170 ;
        RECT 1743.230 1746.990 1744.410 1748.170 ;
        RECT 1741.630 1568.590 1742.810 1569.770 ;
        RECT 1743.230 1568.590 1744.410 1569.770 ;
        RECT 1741.630 1566.990 1742.810 1568.170 ;
        RECT 1743.230 1566.990 1744.410 1568.170 ;
        RECT 1741.630 1388.590 1742.810 1389.770 ;
        RECT 1743.230 1388.590 1744.410 1389.770 ;
        RECT 1741.630 1386.990 1742.810 1388.170 ;
        RECT 1743.230 1386.990 1744.410 1388.170 ;
        RECT 1741.630 1208.590 1742.810 1209.770 ;
        RECT 1743.230 1208.590 1744.410 1209.770 ;
        RECT 1741.630 1206.990 1742.810 1208.170 ;
        RECT 1743.230 1206.990 1744.410 1208.170 ;
        RECT 1741.630 1028.590 1742.810 1029.770 ;
        RECT 1743.230 1028.590 1744.410 1029.770 ;
        RECT 1741.630 1026.990 1742.810 1028.170 ;
        RECT 1743.230 1026.990 1744.410 1028.170 ;
        RECT 1741.630 848.590 1742.810 849.770 ;
        RECT 1743.230 848.590 1744.410 849.770 ;
        RECT 1741.630 846.990 1742.810 848.170 ;
        RECT 1743.230 846.990 1744.410 848.170 ;
        RECT 1741.630 668.590 1742.810 669.770 ;
        RECT 1743.230 668.590 1744.410 669.770 ;
        RECT 1741.630 666.990 1742.810 668.170 ;
        RECT 1743.230 666.990 1744.410 668.170 ;
        RECT 1741.630 488.590 1742.810 489.770 ;
        RECT 1743.230 488.590 1744.410 489.770 ;
        RECT 1741.630 486.990 1742.810 488.170 ;
        RECT 1743.230 486.990 1744.410 488.170 ;
        RECT 1741.630 308.590 1742.810 309.770 ;
        RECT 1743.230 308.590 1744.410 309.770 ;
        RECT 1741.630 306.990 1742.810 308.170 ;
        RECT 1743.230 306.990 1744.410 308.170 ;
        RECT 1741.630 128.590 1742.810 129.770 ;
        RECT 1743.230 128.590 1744.410 129.770 ;
        RECT 1741.630 126.990 1742.810 128.170 ;
        RECT 1743.230 126.990 1744.410 128.170 ;
        RECT 1741.630 -28.460 1742.810 -27.280 ;
        RECT 1743.230 -28.460 1744.410 -27.280 ;
        RECT 1741.630 -30.060 1742.810 -28.880 ;
        RECT 1743.230 -30.060 1744.410 -28.880 ;
        RECT 1921.630 3548.560 1922.810 3549.740 ;
        RECT 1923.230 3548.560 1924.410 3549.740 ;
        RECT 1921.630 3546.960 1922.810 3548.140 ;
        RECT 1923.230 3546.960 1924.410 3548.140 ;
        RECT 1921.630 3368.590 1922.810 3369.770 ;
        RECT 1923.230 3368.590 1924.410 3369.770 ;
        RECT 1921.630 3366.990 1922.810 3368.170 ;
        RECT 1923.230 3366.990 1924.410 3368.170 ;
        RECT 1921.630 3188.590 1922.810 3189.770 ;
        RECT 1923.230 3188.590 1924.410 3189.770 ;
        RECT 1921.630 3186.990 1922.810 3188.170 ;
        RECT 1923.230 3186.990 1924.410 3188.170 ;
        RECT 1921.630 3008.590 1922.810 3009.770 ;
        RECT 1923.230 3008.590 1924.410 3009.770 ;
        RECT 1921.630 3006.990 1922.810 3008.170 ;
        RECT 1923.230 3006.990 1924.410 3008.170 ;
        RECT 1921.630 2828.590 1922.810 2829.770 ;
        RECT 1923.230 2828.590 1924.410 2829.770 ;
        RECT 1921.630 2826.990 1922.810 2828.170 ;
        RECT 1923.230 2826.990 1924.410 2828.170 ;
        RECT 1921.630 2648.590 1922.810 2649.770 ;
        RECT 1923.230 2648.590 1924.410 2649.770 ;
        RECT 1921.630 2646.990 1922.810 2648.170 ;
        RECT 1923.230 2646.990 1924.410 2648.170 ;
        RECT 1921.630 2468.590 1922.810 2469.770 ;
        RECT 1923.230 2468.590 1924.410 2469.770 ;
        RECT 1921.630 2466.990 1922.810 2468.170 ;
        RECT 1923.230 2466.990 1924.410 2468.170 ;
        RECT 1921.630 2288.590 1922.810 2289.770 ;
        RECT 1923.230 2288.590 1924.410 2289.770 ;
        RECT 1921.630 2286.990 1922.810 2288.170 ;
        RECT 1923.230 2286.990 1924.410 2288.170 ;
        RECT 1921.630 2108.590 1922.810 2109.770 ;
        RECT 1923.230 2108.590 1924.410 2109.770 ;
        RECT 1921.630 2106.990 1922.810 2108.170 ;
        RECT 1923.230 2106.990 1924.410 2108.170 ;
        RECT 1921.630 1928.590 1922.810 1929.770 ;
        RECT 1923.230 1928.590 1924.410 1929.770 ;
        RECT 1921.630 1926.990 1922.810 1928.170 ;
        RECT 1923.230 1926.990 1924.410 1928.170 ;
        RECT 1921.630 1748.590 1922.810 1749.770 ;
        RECT 1923.230 1748.590 1924.410 1749.770 ;
        RECT 1921.630 1746.990 1922.810 1748.170 ;
        RECT 1923.230 1746.990 1924.410 1748.170 ;
        RECT 1921.630 1568.590 1922.810 1569.770 ;
        RECT 1923.230 1568.590 1924.410 1569.770 ;
        RECT 1921.630 1566.990 1922.810 1568.170 ;
        RECT 1923.230 1566.990 1924.410 1568.170 ;
        RECT 1921.630 1388.590 1922.810 1389.770 ;
        RECT 1923.230 1388.590 1924.410 1389.770 ;
        RECT 1921.630 1386.990 1922.810 1388.170 ;
        RECT 1923.230 1386.990 1924.410 1388.170 ;
        RECT 1921.630 1208.590 1922.810 1209.770 ;
        RECT 1923.230 1208.590 1924.410 1209.770 ;
        RECT 1921.630 1206.990 1922.810 1208.170 ;
        RECT 1923.230 1206.990 1924.410 1208.170 ;
        RECT 1921.630 1028.590 1922.810 1029.770 ;
        RECT 1923.230 1028.590 1924.410 1029.770 ;
        RECT 1921.630 1026.990 1922.810 1028.170 ;
        RECT 1923.230 1026.990 1924.410 1028.170 ;
        RECT 1921.630 848.590 1922.810 849.770 ;
        RECT 1923.230 848.590 1924.410 849.770 ;
        RECT 1921.630 846.990 1922.810 848.170 ;
        RECT 1923.230 846.990 1924.410 848.170 ;
        RECT 1921.630 668.590 1922.810 669.770 ;
        RECT 1923.230 668.590 1924.410 669.770 ;
        RECT 1921.630 666.990 1922.810 668.170 ;
        RECT 1923.230 666.990 1924.410 668.170 ;
        RECT 1921.630 488.590 1922.810 489.770 ;
        RECT 1923.230 488.590 1924.410 489.770 ;
        RECT 1921.630 486.990 1922.810 488.170 ;
        RECT 1923.230 486.990 1924.410 488.170 ;
        RECT 1921.630 308.590 1922.810 309.770 ;
        RECT 1923.230 308.590 1924.410 309.770 ;
        RECT 1921.630 306.990 1922.810 308.170 ;
        RECT 1923.230 306.990 1924.410 308.170 ;
        RECT 1921.630 128.590 1922.810 129.770 ;
        RECT 1923.230 128.590 1924.410 129.770 ;
        RECT 1921.630 126.990 1922.810 128.170 ;
        RECT 1923.230 126.990 1924.410 128.170 ;
        RECT 1921.630 -28.460 1922.810 -27.280 ;
        RECT 1923.230 -28.460 1924.410 -27.280 ;
        RECT 1921.630 -30.060 1922.810 -28.880 ;
        RECT 1923.230 -30.060 1924.410 -28.880 ;
        RECT 2101.630 3548.560 2102.810 3549.740 ;
        RECT 2103.230 3548.560 2104.410 3549.740 ;
        RECT 2101.630 3546.960 2102.810 3548.140 ;
        RECT 2103.230 3546.960 2104.410 3548.140 ;
        RECT 2101.630 3368.590 2102.810 3369.770 ;
        RECT 2103.230 3368.590 2104.410 3369.770 ;
        RECT 2101.630 3366.990 2102.810 3368.170 ;
        RECT 2103.230 3366.990 2104.410 3368.170 ;
        RECT 2101.630 3188.590 2102.810 3189.770 ;
        RECT 2103.230 3188.590 2104.410 3189.770 ;
        RECT 2101.630 3186.990 2102.810 3188.170 ;
        RECT 2103.230 3186.990 2104.410 3188.170 ;
        RECT 2101.630 3008.590 2102.810 3009.770 ;
        RECT 2103.230 3008.590 2104.410 3009.770 ;
        RECT 2101.630 3006.990 2102.810 3008.170 ;
        RECT 2103.230 3006.990 2104.410 3008.170 ;
        RECT 2101.630 2828.590 2102.810 2829.770 ;
        RECT 2103.230 2828.590 2104.410 2829.770 ;
        RECT 2101.630 2826.990 2102.810 2828.170 ;
        RECT 2103.230 2826.990 2104.410 2828.170 ;
        RECT 2101.630 2648.590 2102.810 2649.770 ;
        RECT 2103.230 2648.590 2104.410 2649.770 ;
        RECT 2101.630 2646.990 2102.810 2648.170 ;
        RECT 2103.230 2646.990 2104.410 2648.170 ;
        RECT 2101.630 2468.590 2102.810 2469.770 ;
        RECT 2103.230 2468.590 2104.410 2469.770 ;
        RECT 2101.630 2466.990 2102.810 2468.170 ;
        RECT 2103.230 2466.990 2104.410 2468.170 ;
        RECT 2101.630 2288.590 2102.810 2289.770 ;
        RECT 2103.230 2288.590 2104.410 2289.770 ;
        RECT 2101.630 2286.990 2102.810 2288.170 ;
        RECT 2103.230 2286.990 2104.410 2288.170 ;
        RECT 2101.630 2108.590 2102.810 2109.770 ;
        RECT 2103.230 2108.590 2104.410 2109.770 ;
        RECT 2101.630 2106.990 2102.810 2108.170 ;
        RECT 2103.230 2106.990 2104.410 2108.170 ;
        RECT 2101.630 1928.590 2102.810 1929.770 ;
        RECT 2103.230 1928.590 2104.410 1929.770 ;
        RECT 2101.630 1926.990 2102.810 1928.170 ;
        RECT 2103.230 1926.990 2104.410 1928.170 ;
        RECT 2101.630 1748.590 2102.810 1749.770 ;
        RECT 2103.230 1748.590 2104.410 1749.770 ;
        RECT 2101.630 1746.990 2102.810 1748.170 ;
        RECT 2103.230 1746.990 2104.410 1748.170 ;
        RECT 2101.630 1568.590 2102.810 1569.770 ;
        RECT 2103.230 1568.590 2104.410 1569.770 ;
        RECT 2101.630 1566.990 2102.810 1568.170 ;
        RECT 2103.230 1566.990 2104.410 1568.170 ;
        RECT 2101.630 1388.590 2102.810 1389.770 ;
        RECT 2103.230 1388.590 2104.410 1389.770 ;
        RECT 2101.630 1386.990 2102.810 1388.170 ;
        RECT 2103.230 1386.990 2104.410 1388.170 ;
        RECT 2101.630 1208.590 2102.810 1209.770 ;
        RECT 2103.230 1208.590 2104.410 1209.770 ;
        RECT 2101.630 1206.990 2102.810 1208.170 ;
        RECT 2103.230 1206.990 2104.410 1208.170 ;
        RECT 2101.630 1028.590 2102.810 1029.770 ;
        RECT 2103.230 1028.590 2104.410 1029.770 ;
        RECT 2101.630 1026.990 2102.810 1028.170 ;
        RECT 2103.230 1026.990 2104.410 1028.170 ;
        RECT 2101.630 848.590 2102.810 849.770 ;
        RECT 2103.230 848.590 2104.410 849.770 ;
        RECT 2101.630 846.990 2102.810 848.170 ;
        RECT 2103.230 846.990 2104.410 848.170 ;
        RECT 2101.630 668.590 2102.810 669.770 ;
        RECT 2103.230 668.590 2104.410 669.770 ;
        RECT 2101.630 666.990 2102.810 668.170 ;
        RECT 2103.230 666.990 2104.410 668.170 ;
        RECT 2101.630 488.590 2102.810 489.770 ;
        RECT 2103.230 488.590 2104.410 489.770 ;
        RECT 2101.630 486.990 2102.810 488.170 ;
        RECT 2103.230 486.990 2104.410 488.170 ;
        RECT 2101.630 308.590 2102.810 309.770 ;
        RECT 2103.230 308.590 2104.410 309.770 ;
        RECT 2101.630 306.990 2102.810 308.170 ;
        RECT 2103.230 306.990 2104.410 308.170 ;
        RECT 2101.630 128.590 2102.810 129.770 ;
        RECT 2103.230 128.590 2104.410 129.770 ;
        RECT 2101.630 126.990 2102.810 128.170 ;
        RECT 2103.230 126.990 2104.410 128.170 ;
        RECT 2101.630 -28.460 2102.810 -27.280 ;
        RECT 2103.230 -28.460 2104.410 -27.280 ;
        RECT 2101.630 -30.060 2102.810 -28.880 ;
        RECT 2103.230 -30.060 2104.410 -28.880 ;
        RECT 2281.630 3548.560 2282.810 3549.740 ;
        RECT 2283.230 3548.560 2284.410 3549.740 ;
        RECT 2281.630 3546.960 2282.810 3548.140 ;
        RECT 2283.230 3546.960 2284.410 3548.140 ;
        RECT 2281.630 3368.590 2282.810 3369.770 ;
        RECT 2283.230 3368.590 2284.410 3369.770 ;
        RECT 2281.630 3366.990 2282.810 3368.170 ;
        RECT 2283.230 3366.990 2284.410 3368.170 ;
        RECT 2281.630 3188.590 2282.810 3189.770 ;
        RECT 2283.230 3188.590 2284.410 3189.770 ;
        RECT 2281.630 3186.990 2282.810 3188.170 ;
        RECT 2283.230 3186.990 2284.410 3188.170 ;
        RECT 2281.630 3008.590 2282.810 3009.770 ;
        RECT 2283.230 3008.590 2284.410 3009.770 ;
        RECT 2281.630 3006.990 2282.810 3008.170 ;
        RECT 2283.230 3006.990 2284.410 3008.170 ;
        RECT 2281.630 2828.590 2282.810 2829.770 ;
        RECT 2283.230 2828.590 2284.410 2829.770 ;
        RECT 2281.630 2826.990 2282.810 2828.170 ;
        RECT 2283.230 2826.990 2284.410 2828.170 ;
        RECT 2281.630 2648.590 2282.810 2649.770 ;
        RECT 2283.230 2648.590 2284.410 2649.770 ;
        RECT 2281.630 2646.990 2282.810 2648.170 ;
        RECT 2283.230 2646.990 2284.410 2648.170 ;
        RECT 2281.630 2468.590 2282.810 2469.770 ;
        RECT 2283.230 2468.590 2284.410 2469.770 ;
        RECT 2281.630 2466.990 2282.810 2468.170 ;
        RECT 2283.230 2466.990 2284.410 2468.170 ;
        RECT 2281.630 2288.590 2282.810 2289.770 ;
        RECT 2283.230 2288.590 2284.410 2289.770 ;
        RECT 2281.630 2286.990 2282.810 2288.170 ;
        RECT 2283.230 2286.990 2284.410 2288.170 ;
        RECT 2281.630 2108.590 2282.810 2109.770 ;
        RECT 2283.230 2108.590 2284.410 2109.770 ;
        RECT 2281.630 2106.990 2282.810 2108.170 ;
        RECT 2283.230 2106.990 2284.410 2108.170 ;
        RECT 2281.630 1928.590 2282.810 1929.770 ;
        RECT 2283.230 1928.590 2284.410 1929.770 ;
        RECT 2281.630 1926.990 2282.810 1928.170 ;
        RECT 2283.230 1926.990 2284.410 1928.170 ;
        RECT 2281.630 1748.590 2282.810 1749.770 ;
        RECT 2283.230 1748.590 2284.410 1749.770 ;
        RECT 2281.630 1746.990 2282.810 1748.170 ;
        RECT 2283.230 1746.990 2284.410 1748.170 ;
        RECT 2281.630 1568.590 2282.810 1569.770 ;
        RECT 2283.230 1568.590 2284.410 1569.770 ;
        RECT 2281.630 1566.990 2282.810 1568.170 ;
        RECT 2283.230 1566.990 2284.410 1568.170 ;
        RECT 2281.630 1388.590 2282.810 1389.770 ;
        RECT 2283.230 1388.590 2284.410 1389.770 ;
        RECT 2281.630 1386.990 2282.810 1388.170 ;
        RECT 2283.230 1386.990 2284.410 1388.170 ;
        RECT 2281.630 1208.590 2282.810 1209.770 ;
        RECT 2283.230 1208.590 2284.410 1209.770 ;
        RECT 2281.630 1206.990 2282.810 1208.170 ;
        RECT 2283.230 1206.990 2284.410 1208.170 ;
        RECT 2281.630 1028.590 2282.810 1029.770 ;
        RECT 2283.230 1028.590 2284.410 1029.770 ;
        RECT 2281.630 1026.990 2282.810 1028.170 ;
        RECT 2283.230 1026.990 2284.410 1028.170 ;
        RECT 2281.630 848.590 2282.810 849.770 ;
        RECT 2283.230 848.590 2284.410 849.770 ;
        RECT 2281.630 846.990 2282.810 848.170 ;
        RECT 2283.230 846.990 2284.410 848.170 ;
        RECT 2281.630 668.590 2282.810 669.770 ;
        RECT 2283.230 668.590 2284.410 669.770 ;
        RECT 2281.630 666.990 2282.810 668.170 ;
        RECT 2283.230 666.990 2284.410 668.170 ;
        RECT 2281.630 488.590 2282.810 489.770 ;
        RECT 2283.230 488.590 2284.410 489.770 ;
        RECT 2281.630 486.990 2282.810 488.170 ;
        RECT 2283.230 486.990 2284.410 488.170 ;
        RECT 2281.630 308.590 2282.810 309.770 ;
        RECT 2283.230 308.590 2284.410 309.770 ;
        RECT 2281.630 306.990 2282.810 308.170 ;
        RECT 2283.230 306.990 2284.410 308.170 ;
        RECT 2281.630 128.590 2282.810 129.770 ;
        RECT 2283.230 128.590 2284.410 129.770 ;
        RECT 2281.630 126.990 2282.810 128.170 ;
        RECT 2283.230 126.990 2284.410 128.170 ;
        RECT 2281.630 -28.460 2282.810 -27.280 ;
        RECT 2283.230 -28.460 2284.410 -27.280 ;
        RECT 2281.630 -30.060 2282.810 -28.880 ;
        RECT 2283.230 -30.060 2284.410 -28.880 ;
        RECT 2461.630 3548.560 2462.810 3549.740 ;
        RECT 2463.230 3548.560 2464.410 3549.740 ;
        RECT 2461.630 3546.960 2462.810 3548.140 ;
        RECT 2463.230 3546.960 2464.410 3548.140 ;
        RECT 2461.630 3368.590 2462.810 3369.770 ;
        RECT 2463.230 3368.590 2464.410 3369.770 ;
        RECT 2461.630 3366.990 2462.810 3368.170 ;
        RECT 2463.230 3366.990 2464.410 3368.170 ;
        RECT 2461.630 3188.590 2462.810 3189.770 ;
        RECT 2463.230 3188.590 2464.410 3189.770 ;
        RECT 2461.630 3186.990 2462.810 3188.170 ;
        RECT 2463.230 3186.990 2464.410 3188.170 ;
        RECT 2461.630 3008.590 2462.810 3009.770 ;
        RECT 2463.230 3008.590 2464.410 3009.770 ;
        RECT 2461.630 3006.990 2462.810 3008.170 ;
        RECT 2463.230 3006.990 2464.410 3008.170 ;
        RECT 2461.630 2828.590 2462.810 2829.770 ;
        RECT 2463.230 2828.590 2464.410 2829.770 ;
        RECT 2461.630 2826.990 2462.810 2828.170 ;
        RECT 2463.230 2826.990 2464.410 2828.170 ;
        RECT 2461.630 2648.590 2462.810 2649.770 ;
        RECT 2463.230 2648.590 2464.410 2649.770 ;
        RECT 2461.630 2646.990 2462.810 2648.170 ;
        RECT 2463.230 2646.990 2464.410 2648.170 ;
        RECT 2461.630 2468.590 2462.810 2469.770 ;
        RECT 2463.230 2468.590 2464.410 2469.770 ;
        RECT 2461.630 2466.990 2462.810 2468.170 ;
        RECT 2463.230 2466.990 2464.410 2468.170 ;
        RECT 2461.630 2288.590 2462.810 2289.770 ;
        RECT 2463.230 2288.590 2464.410 2289.770 ;
        RECT 2461.630 2286.990 2462.810 2288.170 ;
        RECT 2463.230 2286.990 2464.410 2288.170 ;
        RECT 2461.630 2108.590 2462.810 2109.770 ;
        RECT 2463.230 2108.590 2464.410 2109.770 ;
        RECT 2461.630 2106.990 2462.810 2108.170 ;
        RECT 2463.230 2106.990 2464.410 2108.170 ;
        RECT 2461.630 1928.590 2462.810 1929.770 ;
        RECT 2463.230 1928.590 2464.410 1929.770 ;
        RECT 2461.630 1926.990 2462.810 1928.170 ;
        RECT 2463.230 1926.990 2464.410 1928.170 ;
        RECT 2461.630 1748.590 2462.810 1749.770 ;
        RECT 2463.230 1748.590 2464.410 1749.770 ;
        RECT 2461.630 1746.990 2462.810 1748.170 ;
        RECT 2463.230 1746.990 2464.410 1748.170 ;
        RECT 2461.630 1568.590 2462.810 1569.770 ;
        RECT 2463.230 1568.590 2464.410 1569.770 ;
        RECT 2461.630 1566.990 2462.810 1568.170 ;
        RECT 2463.230 1566.990 2464.410 1568.170 ;
        RECT 2461.630 1388.590 2462.810 1389.770 ;
        RECT 2463.230 1388.590 2464.410 1389.770 ;
        RECT 2461.630 1386.990 2462.810 1388.170 ;
        RECT 2463.230 1386.990 2464.410 1388.170 ;
        RECT 2461.630 1208.590 2462.810 1209.770 ;
        RECT 2463.230 1208.590 2464.410 1209.770 ;
        RECT 2461.630 1206.990 2462.810 1208.170 ;
        RECT 2463.230 1206.990 2464.410 1208.170 ;
        RECT 2461.630 1028.590 2462.810 1029.770 ;
        RECT 2463.230 1028.590 2464.410 1029.770 ;
        RECT 2461.630 1026.990 2462.810 1028.170 ;
        RECT 2463.230 1026.990 2464.410 1028.170 ;
        RECT 2461.630 848.590 2462.810 849.770 ;
        RECT 2463.230 848.590 2464.410 849.770 ;
        RECT 2461.630 846.990 2462.810 848.170 ;
        RECT 2463.230 846.990 2464.410 848.170 ;
        RECT 2461.630 668.590 2462.810 669.770 ;
        RECT 2463.230 668.590 2464.410 669.770 ;
        RECT 2461.630 666.990 2462.810 668.170 ;
        RECT 2463.230 666.990 2464.410 668.170 ;
        RECT 2461.630 488.590 2462.810 489.770 ;
        RECT 2463.230 488.590 2464.410 489.770 ;
        RECT 2461.630 486.990 2462.810 488.170 ;
        RECT 2463.230 486.990 2464.410 488.170 ;
        RECT 2461.630 308.590 2462.810 309.770 ;
        RECT 2463.230 308.590 2464.410 309.770 ;
        RECT 2461.630 306.990 2462.810 308.170 ;
        RECT 2463.230 306.990 2464.410 308.170 ;
        RECT 2461.630 128.590 2462.810 129.770 ;
        RECT 2463.230 128.590 2464.410 129.770 ;
        RECT 2461.630 126.990 2462.810 128.170 ;
        RECT 2463.230 126.990 2464.410 128.170 ;
        RECT 2461.630 -28.460 2462.810 -27.280 ;
        RECT 2463.230 -28.460 2464.410 -27.280 ;
        RECT 2461.630 -30.060 2462.810 -28.880 ;
        RECT 2463.230 -30.060 2464.410 -28.880 ;
        RECT 2641.630 3548.560 2642.810 3549.740 ;
        RECT 2643.230 3548.560 2644.410 3549.740 ;
        RECT 2641.630 3546.960 2642.810 3548.140 ;
        RECT 2643.230 3546.960 2644.410 3548.140 ;
        RECT 2641.630 3368.590 2642.810 3369.770 ;
        RECT 2643.230 3368.590 2644.410 3369.770 ;
        RECT 2641.630 3366.990 2642.810 3368.170 ;
        RECT 2643.230 3366.990 2644.410 3368.170 ;
        RECT 2641.630 3188.590 2642.810 3189.770 ;
        RECT 2643.230 3188.590 2644.410 3189.770 ;
        RECT 2641.630 3186.990 2642.810 3188.170 ;
        RECT 2643.230 3186.990 2644.410 3188.170 ;
        RECT 2641.630 3008.590 2642.810 3009.770 ;
        RECT 2643.230 3008.590 2644.410 3009.770 ;
        RECT 2641.630 3006.990 2642.810 3008.170 ;
        RECT 2643.230 3006.990 2644.410 3008.170 ;
        RECT 2641.630 2828.590 2642.810 2829.770 ;
        RECT 2643.230 2828.590 2644.410 2829.770 ;
        RECT 2641.630 2826.990 2642.810 2828.170 ;
        RECT 2643.230 2826.990 2644.410 2828.170 ;
        RECT 2641.630 2648.590 2642.810 2649.770 ;
        RECT 2643.230 2648.590 2644.410 2649.770 ;
        RECT 2641.630 2646.990 2642.810 2648.170 ;
        RECT 2643.230 2646.990 2644.410 2648.170 ;
        RECT 2641.630 2468.590 2642.810 2469.770 ;
        RECT 2643.230 2468.590 2644.410 2469.770 ;
        RECT 2641.630 2466.990 2642.810 2468.170 ;
        RECT 2643.230 2466.990 2644.410 2468.170 ;
        RECT 2641.630 2288.590 2642.810 2289.770 ;
        RECT 2643.230 2288.590 2644.410 2289.770 ;
        RECT 2641.630 2286.990 2642.810 2288.170 ;
        RECT 2643.230 2286.990 2644.410 2288.170 ;
        RECT 2641.630 2108.590 2642.810 2109.770 ;
        RECT 2643.230 2108.590 2644.410 2109.770 ;
        RECT 2641.630 2106.990 2642.810 2108.170 ;
        RECT 2643.230 2106.990 2644.410 2108.170 ;
        RECT 2641.630 1928.590 2642.810 1929.770 ;
        RECT 2643.230 1928.590 2644.410 1929.770 ;
        RECT 2641.630 1926.990 2642.810 1928.170 ;
        RECT 2643.230 1926.990 2644.410 1928.170 ;
        RECT 2641.630 1748.590 2642.810 1749.770 ;
        RECT 2643.230 1748.590 2644.410 1749.770 ;
        RECT 2641.630 1746.990 2642.810 1748.170 ;
        RECT 2643.230 1746.990 2644.410 1748.170 ;
        RECT 2641.630 1568.590 2642.810 1569.770 ;
        RECT 2643.230 1568.590 2644.410 1569.770 ;
        RECT 2641.630 1566.990 2642.810 1568.170 ;
        RECT 2643.230 1566.990 2644.410 1568.170 ;
        RECT 2641.630 1388.590 2642.810 1389.770 ;
        RECT 2643.230 1388.590 2644.410 1389.770 ;
        RECT 2641.630 1386.990 2642.810 1388.170 ;
        RECT 2643.230 1386.990 2644.410 1388.170 ;
        RECT 2641.630 1208.590 2642.810 1209.770 ;
        RECT 2643.230 1208.590 2644.410 1209.770 ;
        RECT 2641.630 1206.990 2642.810 1208.170 ;
        RECT 2643.230 1206.990 2644.410 1208.170 ;
        RECT 2641.630 1028.590 2642.810 1029.770 ;
        RECT 2643.230 1028.590 2644.410 1029.770 ;
        RECT 2641.630 1026.990 2642.810 1028.170 ;
        RECT 2643.230 1026.990 2644.410 1028.170 ;
        RECT 2641.630 848.590 2642.810 849.770 ;
        RECT 2643.230 848.590 2644.410 849.770 ;
        RECT 2641.630 846.990 2642.810 848.170 ;
        RECT 2643.230 846.990 2644.410 848.170 ;
        RECT 2641.630 668.590 2642.810 669.770 ;
        RECT 2643.230 668.590 2644.410 669.770 ;
        RECT 2641.630 666.990 2642.810 668.170 ;
        RECT 2643.230 666.990 2644.410 668.170 ;
        RECT 2641.630 488.590 2642.810 489.770 ;
        RECT 2643.230 488.590 2644.410 489.770 ;
        RECT 2641.630 486.990 2642.810 488.170 ;
        RECT 2643.230 486.990 2644.410 488.170 ;
        RECT 2641.630 308.590 2642.810 309.770 ;
        RECT 2643.230 308.590 2644.410 309.770 ;
        RECT 2641.630 306.990 2642.810 308.170 ;
        RECT 2643.230 306.990 2644.410 308.170 ;
        RECT 2641.630 128.590 2642.810 129.770 ;
        RECT 2643.230 128.590 2644.410 129.770 ;
        RECT 2641.630 126.990 2642.810 128.170 ;
        RECT 2643.230 126.990 2644.410 128.170 ;
        RECT 2641.630 -28.460 2642.810 -27.280 ;
        RECT 2643.230 -28.460 2644.410 -27.280 ;
        RECT 2641.630 -30.060 2642.810 -28.880 ;
        RECT 2643.230 -30.060 2644.410 -28.880 ;
        RECT 2821.630 3548.560 2822.810 3549.740 ;
        RECT 2823.230 3548.560 2824.410 3549.740 ;
        RECT 2821.630 3546.960 2822.810 3548.140 ;
        RECT 2823.230 3546.960 2824.410 3548.140 ;
        RECT 2821.630 3368.590 2822.810 3369.770 ;
        RECT 2823.230 3368.590 2824.410 3369.770 ;
        RECT 2821.630 3366.990 2822.810 3368.170 ;
        RECT 2823.230 3366.990 2824.410 3368.170 ;
        RECT 2821.630 3188.590 2822.810 3189.770 ;
        RECT 2823.230 3188.590 2824.410 3189.770 ;
        RECT 2821.630 3186.990 2822.810 3188.170 ;
        RECT 2823.230 3186.990 2824.410 3188.170 ;
        RECT 2821.630 3008.590 2822.810 3009.770 ;
        RECT 2823.230 3008.590 2824.410 3009.770 ;
        RECT 2821.630 3006.990 2822.810 3008.170 ;
        RECT 2823.230 3006.990 2824.410 3008.170 ;
        RECT 2821.630 2828.590 2822.810 2829.770 ;
        RECT 2823.230 2828.590 2824.410 2829.770 ;
        RECT 2821.630 2826.990 2822.810 2828.170 ;
        RECT 2823.230 2826.990 2824.410 2828.170 ;
        RECT 2821.630 2648.590 2822.810 2649.770 ;
        RECT 2823.230 2648.590 2824.410 2649.770 ;
        RECT 2821.630 2646.990 2822.810 2648.170 ;
        RECT 2823.230 2646.990 2824.410 2648.170 ;
        RECT 2821.630 2468.590 2822.810 2469.770 ;
        RECT 2823.230 2468.590 2824.410 2469.770 ;
        RECT 2821.630 2466.990 2822.810 2468.170 ;
        RECT 2823.230 2466.990 2824.410 2468.170 ;
        RECT 2821.630 2288.590 2822.810 2289.770 ;
        RECT 2823.230 2288.590 2824.410 2289.770 ;
        RECT 2821.630 2286.990 2822.810 2288.170 ;
        RECT 2823.230 2286.990 2824.410 2288.170 ;
        RECT 2821.630 2108.590 2822.810 2109.770 ;
        RECT 2823.230 2108.590 2824.410 2109.770 ;
        RECT 2821.630 2106.990 2822.810 2108.170 ;
        RECT 2823.230 2106.990 2824.410 2108.170 ;
        RECT 2821.630 1928.590 2822.810 1929.770 ;
        RECT 2823.230 1928.590 2824.410 1929.770 ;
        RECT 2821.630 1926.990 2822.810 1928.170 ;
        RECT 2823.230 1926.990 2824.410 1928.170 ;
        RECT 2821.630 1748.590 2822.810 1749.770 ;
        RECT 2823.230 1748.590 2824.410 1749.770 ;
        RECT 2821.630 1746.990 2822.810 1748.170 ;
        RECT 2823.230 1746.990 2824.410 1748.170 ;
        RECT 2821.630 1568.590 2822.810 1569.770 ;
        RECT 2823.230 1568.590 2824.410 1569.770 ;
        RECT 2821.630 1566.990 2822.810 1568.170 ;
        RECT 2823.230 1566.990 2824.410 1568.170 ;
        RECT 2821.630 1388.590 2822.810 1389.770 ;
        RECT 2823.230 1388.590 2824.410 1389.770 ;
        RECT 2821.630 1386.990 2822.810 1388.170 ;
        RECT 2823.230 1386.990 2824.410 1388.170 ;
        RECT 2821.630 1208.590 2822.810 1209.770 ;
        RECT 2823.230 1208.590 2824.410 1209.770 ;
        RECT 2821.630 1206.990 2822.810 1208.170 ;
        RECT 2823.230 1206.990 2824.410 1208.170 ;
        RECT 2821.630 1028.590 2822.810 1029.770 ;
        RECT 2823.230 1028.590 2824.410 1029.770 ;
        RECT 2821.630 1026.990 2822.810 1028.170 ;
        RECT 2823.230 1026.990 2824.410 1028.170 ;
        RECT 2821.630 848.590 2822.810 849.770 ;
        RECT 2823.230 848.590 2824.410 849.770 ;
        RECT 2821.630 846.990 2822.810 848.170 ;
        RECT 2823.230 846.990 2824.410 848.170 ;
        RECT 2821.630 668.590 2822.810 669.770 ;
        RECT 2823.230 668.590 2824.410 669.770 ;
        RECT 2821.630 666.990 2822.810 668.170 ;
        RECT 2823.230 666.990 2824.410 668.170 ;
        RECT 2821.630 488.590 2822.810 489.770 ;
        RECT 2823.230 488.590 2824.410 489.770 ;
        RECT 2821.630 486.990 2822.810 488.170 ;
        RECT 2823.230 486.990 2824.410 488.170 ;
        RECT 2821.630 308.590 2822.810 309.770 ;
        RECT 2823.230 308.590 2824.410 309.770 ;
        RECT 2821.630 306.990 2822.810 308.170 ;
        RECT 2823.230 306.990 2824.410 308.170 ;
        RECT 2821.630 128.590 2822.810 129.770 ;
        RECT 2823.230 128.590 2824.410 129.770 ;
        RECT 2821.630 126.990 2822.810 128.170 ;
        RECT 2823.230 126.990 2824.410 128.170 ;
        RECT 2821.630 -28.460 2822.810 -27.280 ;
        RECT 2823.230 -28.460 2824.410 -27.280 ;
        RECT 2821.630 -30.060 2822.810 -28.880 ;
        RECT 2823.230 -30.060 2824.410 -28.880 ;
        RECT 2952.260 3548.560 2953.440 3549.740 ;
        RECT 2953.860 3548.560 2955.040 3549.740 ;
        RECT 2952.260 3546.960 2953.440 3548.140 ;
        RECT 2953.860 3546.960 2955.040 3548.140 ;
        RECT 2952.260 3368.590 2953.440 3369.770 ;
        RECT 2953.860 3368.590 2955.040 3369.770 ;
        RECT 2952.260 3366.990 2953.440 3368.170 ;
        RECT 2953.860 3366.990 2955.040 3368.170 ;
        RECT 2952.260 3188.590 2953.440 3189.770 ;
        RECT 2953.860 3188.590 2955.040 3189.770 ;
        RECT 2952.260 3186.990 2953.440 3188.170 ;
        RECT 2953.860 3186.990 2955.040 3188.170 ;
        RECT 2952.260 3008.590 2953.440 3009.770 ;
        RECT 2953.860 3008.590 2955.040 3009.770 ;
        RECT 2952.260 3006.990 2953.440 3008.170 ;
        RECT 2953.860 3006.990 2955.040 3008.170 ;
        RECT 2952.260 2828.590 2953.440 2829.770 ;
        RECT 2953.860 2828.590 2955.040 2829.770 ;
        RECT 2952.260 2826.990 2953.440 2828.170 ;
        RECT 2953.860 2826.990 2955.040 2828.170 ;
        RECT 2952.260 2648.590 2953.440 2649.770 ;
        RECT 2953.860 2648.590 2955.040 2649.770 ;
        RECT 2952.260 2646.990 2953.440 2648.170 ;
        RECT 2953.860 2646.990 2955.040 2648.170 ;
        RECT 2952.260 2468.590 2953.440 2469.770 ;
        RECT 2953.860 2468.590 2955.040 2469.770 ;
        RECT 2952.260 2466.990 2953.440 2468.170 ;
        RECT 2953.860 2466.990 2955.040 2468.170 ;
        RECT 2952.260 2288.590 2953.440 2289.770 ;
        RECT 2953.860 2288.590 2955.040 2289.770 ;
        RECT 2952.260 2286.990 2953.440 2288.170 ;
        RECT 2953.860 2286.990 2955.040 2288.170 ;
        RECT 2952.260 2108.590 2953.440 2109.770 ;
        RECT 2953.860 2108.590 2955.040 2109.770 ;
        RECT 2952.260 2106.990 2953.440 2108.170 ;
        RECT 2953.860 2106.990 2955.040 2108.170 ;
        RECT 2952.260 1928.590 2953.440 1929.770 ;
        RECT 2953.860 1928.590 2955.040 1929.770 ;
        RECT 2952.260 1926.990 2953.440 1928.170 ;
        RECT 2953.860 1926.990 2955.040 1928.170 ;
        RECT 2952.260 1748.590 2953.440 1749.770 ;
        RECT 2953.860 1748.590 2955.040 1749.770 ;
        RECT 2952.260 1746.990 2953.440 1748.170 ;
        RECT 2953.860 1746.990 2955.040 1748.170 ;
        RECT 2952.260 1568.590 2953.440 1569.770 ;
        RECT 2953.860 1568.590 2955.040 1569.770 ;
        RECT 2952.260 1566.990 2953.440 1568.170 ;
        RECT 2953.860 1566.990 2955.040 1568.170 ;
        RECT 2952.260 1388.590 2953.440 1389.770 ;
        RECT 2953.860 1388.590 2955.040 1389.770 ;
        RECT 2952.260 1386.990 2953.440 1388.170 ;
        RECT 2953.860 1386.990 2955.040 1388.170 ;
        RECT 2952.260 1208.590 2953.440 1209.770 ;
        RECT 2953.860 1208.590 2955.040 1209.770 ;
        RECT 2952.260 1206.990 2953.440 1208.170 ;
        RECT 2953.860 1206.990 2955.040 1208.170 ;
        RECT 2952.260 1028.590 2953.440 1029.770 ;
        RECT 2953.860 1028.590 2955.040 1029.770 ;
        RECT 2952.260 1026.990 2953.440 1028.170 ;
        RECT 2953.860 1026.990 2955.040 1028.170 ;
        RECT 2952.260 848.590 2953.440 849.770 ;
        RECT 2953.860 848.590 2955.040 849.770 ;
        RECT 2952.260 846.990 2953.440 848.170 ;
        RECT 2953.860 846.990 2955.040 848.170 ;
        RECT 2952.260 668.590 2953.440 669.770 ;
        RECT 2953.860 668.590 2955.040 669.770 ;
        RECT 2952.260 666.990 2953.440 668.170 ;
        RECT 2953.860 666.990 2955.040 668.170 ;
        RECT 2952.260 488.590 2953.440 489.770 ;
        RECT 2953.860 488.590 2955.040 489.770 ;
        RECT 2952.260 486.990 2953.440 488.170 ;
        RECT 2953.860 486.990 2955.040 488.170 ;
        RECT 2952.260 308.590 2953.440 309.770 ;
        RECT 2953.860 308.590 2955.040 309.770 ;
        RECT 2952.260 306.990 2953.440 308.170 ;
        RECT 2953.860 306.990 2955.040 308.170 ;
        RECT 2952.260 128.590 2953.440 129.770 ;
        RECT 2953.860 128.590 2955.040 129.770 ;
        RECT 2952.260 126.990 2953.440 128.170 ;
        RECT 2953.860 126.990 2955.040 128.170 ;
        RECT 2952.260 -28.460 2953.440 -27.280 ;
        RECT 2953.860 -28.460 2955.040 -27.280 ;
        RECT 2952.260 -30.060 2953.440 -28.880 ;
        RECT 2953.860 -30.060 2955.040 -28.880 ;
      LAYER met5 ;
        RECT -35.580 3546.800 2955.200 3549.900 ;
        RECT -45.180 3366.830 2964.800 3369.930 ;
        RECT -45.180 3186.830 2964.800 3189.930 ;
        RECT -45.180 3006.830 2964.800 3009.930 ;
        RECT -45.180 2826.830 2964.800 2829.930 ;
        RECT -45.180 2646.830 2964.800 2649.930 ;
        RECT -45.180 2466.830 2964.800 2469.930 ;
        RECT -45.180 2286.830 2964.800 2289.930 ;
        RECT -45.180 2106.830 2964.800 2109.930 ;
        RECT -45.180 1926.830 2964.800 1929.930 ;
        RECT -45.180 1746.830 2964.800 1749.930 ;
        RECT -45.180 1566.830 2964.800 1569.930 ;
        RECT -45.180 1386.830 2964.800 1389.930 ;
        RECT -45.180 1206.830 2964.800 1209.930 ;
        RECT -45.180 1026.830 2964.800 1029.930 ;
        RECT -45.180 846.830 2964.800 849.930 ;
        RECT -45.180 666.830 2964.800 669.930 ;
        RECT -45.180 486.830 2964.800 489.930 ;
        RECT -45.180 306.830 2964.800 309.930 ;
        RECT -45.180 126.830 2964.800 129.930 ;
        RECT -35.580 -30.220 2955.200 -27.120 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -45.180 -39.820 -42.080 3559.500 ;
        RECT 166.470 -39.820 169.570 3559.500 ;
        RECT 346.470 -39.820 349.570 3559.500 ;
        RECT 526.470 760.000 529.570 3559.500 ;
        RECT 526.470 -39.820 529.570 490.000 ;
        RECT 706.470 -39.820 709.570 3559.500 ;
        RECT 886.470 -39.820 889.570 3559.500 ;
        RECT 1066.470 -39.820 1069.570 3559.500 ;
        RECT 1246.470 -39.820 1249.570 3559.500 ;
        RECT 1426.470 -39.820 1429.570 3559.500 ;
        RECT 1606.470 -39.820 1609.570 3559.500 ;
        RECT 1786.470 -39.820 1789.570 3559.500 ;
        RECT 1966.470 -39.820 1969.570 3559.500 ;
        RECT 2146.470 -39.820 2149.570 3559.500 ;
        RECT 2326.470 -39.820 2329.570 3559.500 ;
        RECT 2506.470 -39.820 2509.570 3559.500 ;
        RECT 2686.470 -39.820 2689.570 3559.500 ;
        RECT 2866.470 -39.820 2869.570 3559.500 ;
        RECT 2961.700 -39.820 2964.800 3559.500 ;
      LAYER via4 ;
        RECT -45.020 3558.160 -43.840 3559.340 ;
        RECT -43.420 3558.160 -42.240 3559.340 ;
        RECT -45.020 3556.560 -43.840 3557.740 ;
        RECT -43.420 3556.560 -42.240 3557.740 ;
        RECT -45.020 3413.590 -43.840 3414.770 ;
        RECT -43.420 3413.590 -42.240 3414.770 ;
        RECT -45.020 3411.990 -43.840 3413.170 ;
        RECT -43.420 3411.990 -42.240 3413.170 ;
        RECT -45.020 3233.590 -43.840 3234.770 ;
        RECT -43.420 3233.590 -42.240 3234.770 ;
        RECT -45.020 3231.990 -43.840 3233.170 ;
        RECT -43.420 3231.990 -42.240 3233.170 ;
        RECT -45.020 3053.590 -43.840 3054.770 ;
        RECT -43.420 3053.590 -42.240 3054.770 ;
        RECT -45.020 3051.990 -43.840 3053.170 ;
        RECT -43.420 3051.990 -42.240 3053.170 ;
        RECT -45.020 2873.590 -43.840 2874.770 ;
        RECT -43.420 2873.590 -42.240 2874.770 ;
        RECT -45.020 2871.990 -43.840 2873.170 ;
        RECT -43.420 2871.990 -42.240 2873.170 ;
        RECT -45.020 2693.590 -43.840 2694.770 ;
        RECT -43.420 2693.590 -42.240 2694.770 ;
        RECT -45.020 2691.990 -43.840 2693.170 ;
        RECT -43.420 2691.990 -42.240 2693.170 ;
        RECT -45.020 2513.590 -43.840 2514.770 ;
        RECT -43.420 2513.590 -42.240 2514.770 ;
        RECT -45.020 2511.990 -43.840 2513.170 ;
        RECT -43.420 2511.990 -42.240 2513.170 ;
        RECT -45.020 2333.590 -43.840 2334.770 ;
        RECT -43.420 2333.590 -42.240 2334.770 ;
        RECT -45.020 2331.990 -43.840 2333.170 ;
        RECT -43.420 2331.990 -42.240 2333.170 ;
        RECT -45.020 2153.590 -43.840 2154.770 ;
        RECT -43.420 2153.590 -42.240 2154.770 ;
        RECT -45.020 2151.990 -43.840 2153.170 ;
        RECT -43.420 2151.990 -42.240 2153.170 ;
        RECT -45.020 1973.590 -43.840 1974.770 ;
        RECT -43.420 1973.590 -42.240 1974.770 ;
        RECT -45.020 1971.990 -43.840 1973.170 ;
        RECT -43.420 1971.990 -42.240 1973.170 ;
        RECT -45.020 1793.590 -43.840 1794.770 ;
        RECT -43.420 1793.590 -42.240 1794.770 ;
        RECT -45.020 1791.990 -43.840 1793.170 ;
        RECT -43.420 1791.990 -42.240 1793.170 ;
        RECT -45.020 1613.590 -43.840 1614.770 ;
        RECT -43.420 1613.590 -42.240 1614.770 ;
        RECT -45.020 1611.990 -43.840 1613.170 ;
        RECT -43.420 1611.990 -42.240 1613.170 ;
        RECT -45.020 1433.590 -43.840 1434.770 ;
        RECT -43.420 1433.590 -42.240 1434.770 ;
        RECT -45.020 1431.990 -43.840 1433.170 ;
        RECT -43.420 1431.990 -42.240 1433.170 ;
        RECT -45.020 1253.590 -43.840 1254.770 ;
        RECT -43.420 1253.590 -42.240 1254.770 ;
        RECT -45.020 1251.990 -43.840 1253.170 ;
        RECT -43.420 1251.990 -42.240 1253.170 ;
        RECT -45.020 1073.590 -43.840 1074.770 ;
        RECT -43.420 1073.590 -42.240 1074.770 ;
        RECT -45.020 1071.990 -43.840 1073.170 ;
        RECT -43.420 1071.990 -42.240 1073.170 ;
        RECT -45.020 893.590 -43.840 894.770 ;
        RECT -43.420 893.590 -42.240 894.770 ;
        RECT -45.020 891.990 -43.840 893.170 ;
        RECT -43.420 891.990 -42.240 893.170 ;
        RECT -45.020 713.590 -43.840 714.770 ;
        RECT -43.420 713.590 -42.240 714.770 ;
        RECT -45.020 711.990 -43.840 713.170 ;
        RECT -43.420 711.990 -42.240 713.170 ;
        RECT -45.020 533.590 -43.840 534.770 ;
        RECT -43.420 533.590 -42.240 534.770 ;
        RECT -45.020 531.990 -43.840 533.170 ;
        RECT -43.420 531.990 -42.240 533.170 ;
        RECT -45.020 353.590 -43.840 354.770 ;
        RECT -43.420 353.590 -42.240 354.770 ;
        RECT -45.020 351.990 -43.840 353.170 ;
        RECT -43.420 351.990 -42.240 353.170 ;
        RECT -45.020 173.590 -43.840 174.770 ;
        RECT -43.420 173.590 -42.240 174.770 ;
        RECT -45.020 171.990 -43.840 173.170 ;
        RECT -43.420 171.990 -42.240 173.170 ;
        RECT -45.020 -38.060 -43.840 -36.880 ;
        RECT -43.420 -38.060 -42.240 -36.880 ;
        RECT -45.020 -39.660 -43.840 -38.480 ;
        RECT -43.420 -39.660 -42.240 -38.480 ;
        RECT 166.630 3558.160 167.810 3559.340 ;
        RECT 168.230 3558.160 169.410 3559.340 ;
        RECT 166.630 3556.560 167.810 3557.740 ;
        RECT 168.230 3556.560 169.410 3557.740 ;
        RECT 166.630 3413.590 167.810 3414.770 ;
        RECT 168.230 3413.590 169.410 3414.770 ;
        RECT 166.630 3411.990 167.810 3413.170 ;
        RECT 168.230 3411.990 169.410 3413.170 ;
        RECT 166.630 3233.590 167.810 3234.770 ;
        RECT 168.230 3233.590 169.410 3234.770 ;
        RECT 166.630 3231.990 167.810 3233.170 ;
        RECT 168.230 3231.990 169.410 3233.170 ;
        RECT 166.630 3053.590 167.810 3054.770 ;
        RECT 168.230 3053.590 169.410 3054.770 ;
        RECT 166.630 3051.990 167.810 3053.170 ;
        RECT 168.230 3051.990 169.410 3053.170 ;
        RECT 166.630 2873.590 167.810 2874.770 ;
        RECT 168.230 2873.590 169.410 2874.770 ;
        RECT 166.630 2871.990 167.810 2873.170 ;
        RECT 168.230 2871.990 169.410 2873.170 ;
        RECT 166.630 2693.590 167.810 2694.770 ;
        RECT 168.230 2693.590 169.410 2694.770 ;
        RECT 166.630 2691.990 167.810 2693.170 ;
        RECT 168.230 2691.990 169.410 2693.170 ;
        RECT 166.630 2513.590 167.810 2514.770 ;
        RECT 168.230 2513.590 169.410 2514.770 ;
        RECT 166.630 2511.990 167.810 2513.170 ;
        RECT 168.230 2511.990 169.410 2513.170 ;
        RECT 166.630 2333.590 167.810 2334.770 ;
        RECT 168.230 2333.590 169.410 2334.770 ;
        RECT 166.630 2331.990 167.810 2333.170 ;
        RECT 168.230 2331.990 169.410 2333.170 ;
        RECT 166.630 2153.590 167.810 2154.770 ;
        RECT 168.230 2153.590 169.410 2154.770 ;
        RECT 166.630 2151.990 167.810 2153.170 ;
        RECT 168.230 2151.990 169.410 2153.170 ;
        RECT 166.630 1973.590 167.810 1974.770 ;
        RECT 168.230 1973.590 169.410 1974.770 ;
        RECT 166.630 1971.990 167.810 1973.170 ;
        RECT 168.230 1971.990 169.410 1973.170 ;
        RECT 166.630 1793.590 167.810 1794.770 ;
        RECT 168.230 1793.590 169.410 1794.770 ;
        RECT 166.630 1791.990 167.810 1793.170 ;
        RECT 168.230 1791.990 169.410 1793.170 ;
        RECT 166.630 1613.590 167.810 1614.770 ;
        RECT 168.230 1613.590 169.410 1614.770 ;
        RECT 166.630 1611.990 167.810 1613.170 ;
        RECT 168.230 1611.990 169.410 1613.170 ;
        RECT 166.630 1433.590 167.810 1434.770 ;
        RECT 168.230 1433.590 169.410 1434.770 ;
        RECT 166.630 1431.990 167.810 1433.170 ;
        RECT 168.230 1431.990 169.410 1433.170 ;
        RECT 166.630 1253.590 167.810 1254.770 ;
        RECT 168.230 1253.590 169.410 1254.770 ;
        RECT 166.630 1251.990 167.810 1253.170 ;
        RECT 168.230 1251.990 169.410 1253.170 ;
        RECT 166.630 1073.590 167.810 1074.770 ;
        RECT 168.230 1073.590 169.410 1074.770 ;
        RECT 166.630 1071.990 167.810 1073.170 ;
        RECT 168.230 1071.990 169.410 1073.170 ;
        RECT 166.630 893.590 167.810 894.770 ;
        RECT 168.230 893.590 169.410 894.770 ;
        RECT 166.630 891.990 167.810 893.170 ;
        RECT 168.230 891.990 169.410 893.170 ;
        RECT 166.630 713.590 167.810 714.770 ;
        RECT 168.230 713.590 169.410 714.770 ;
        RECT 166.630 711.990 167.810 713.170 ;
        RECT 168.230 711.990 169.410 713.170 ;
        RECT 166.630 533.590 167.810 534.770 ;
        RECT 168.230 533.590 169.410 534.770 ;
        RECT 166.630 531.990 167.810 533.170 ;
        RECT 168.230 531.990 169.410 533.170 ;
        RECT 166.630 353.590 167.810 354.770 ;
        RECT 168.230 353.590 169.410 354.770 ;
        RECT 166.630 351.990 167.810 353.170 ;
        RECT 168.230 351.990 169.410 353.170 ;
        RECT 166.630 173.590 167.810 174.770 ;
        RECT 168.230 173.590 169.410 174.770 ;
        RECT 166.630 171.990 167.810 173.170 ;
        RECT 168.230 171.990 169.410 173.170 ;
        RECT 166.630 -38.060 167.810 -36.880 ;
        RECT 168.230 -38.060 169.410 -36.880 ;
        RECT 166.630 -39.660 167.810 -38.480 ;
        RECT 168.230 -39.660 169.410 -38.480 ;
        RECT 346.630 3558.160 347.810 3559.340 ;
        RECT 348.230 3558.160 349.410 3559.340 ;
        RECT 346.630 3556.560 347.810 3557.740 ;
        RECT 348.230 3556.560 349.410 3557.740 ;
        RECT 346.630 3413.590 347.810 3414.770 ;
        RECT 348.230 3413.590 349.410 3414.770 ;
        RECT 346.630 3411.990 347.810 3413.170 ;
        RECT 348.230 3411.990 349.410 3413.170 ;
        RECT 346.630 3233.590 347.810 3234.770 ;
        RECT 348.230 3233.590 349.410 3234.770 ;
        RECT 346.630 3231.990 347.810 3233.170 ;
        RECT 348.230 3231.990 349.410 3233.170 ;
        RECT 346.630 3053.590 347.810 3054.770 ;
        RECT 348.230 3053.590 349.410 3054.770 ;
        RECT 346.630 3051.990 347.810 3053.170 ;
        RECT 348.230 3051.990 349.410 3053.170 ;
        RECT 346.630 2873.590 347.810 2874.770 ;
        RECT 348.230 2873.590 349.410 2874.770 ;
        RECT 346.630 2871.990 347.810 2873.170 ;
        RECT 348.230 2871.990 349.410 2873.170 ;
        RECT 346.630 2693.590 347.810 2694.770 ;
        RECT 348.230 2693.590 349.410 2694.770 ;
        RECT 346.630 2691.990 347.810 2693.170 ;
        RECT 348.230 2691.990 349.410 2693.170 ;
        RECT 346.630 2513.590 347.810 2514.770 ;
        RECT 348.230 2513.590 349.410 2514.770 ;
        RECT 346.630 2511.990 347.810 2513.170 ;
        RECT 348.230 2511.990 349.410 2513.170 ;
        RECT 346.630 2333.590 347.810 2334.770 ;
        RECT 348.230 2333.590 349.410 2334.770 ;
        RECT 346.630 2331.990 347.810 2333.170 ;
        RECT 348.230 2331.990 349.410 2333.170 ;
        RECT 346.630 2153.590 347.810 2154.770 ;
        RECT 348.230 2153.590 349.410 2154.770 ;
        RECT 346.630 2151.990 347.810 2153.170 ;
        RECT 348.230 2151.990 349.410 2153.170 ;
        RECT 346.630 1973.590 347.810 1974.770 ;
        RECT 348.230 1973.590 349.410 1974.770 ;
        RECT 346.630 1971.990 347.810 1973.170 ;
        RECT 348.230 1971.990 349.410 1973.170 ;
        RECT 346.630 1793.590 347.810 1794.770 ;
        RECT 348.230 1793.590 349.410 1794.770 ;
        RECT 346.630 1791.990 347.810 1793.170 ;
        RECT 348.230 1791.990 349.410 1793.170 ;
        RECT 346.630 1613.590 347.810 1614.770 ;
        RECT 348.230 1613.590 349.410 1614.770 ;
        RECT 346.630 1611.990 347.810 1613.170 ;
        RECT 348.230 1611.990 349.410 1613.170 ;
        RECT 346.630 1433.590 347.810 1434.770 ;
        RECT 348.230 1433.590 349.410 1434.770 ;
        RECT 346.630 1431.990 347.810 1433.170 ;
        RECT 348.230 1431.990 349.410 1433.170 ;
        RECT 346.630 1253.590 347.810 1254.770 ;
        RECT 348.230 1253.590 349.410 1254.770 ;
        RECT 346.630 1251.990 347.810 1253.170 ;
        RECT 348.230 1251.990 349.410 1253.170 ;
        RECT 346.630 1073.590 347.810 1074.770 ;
        RECT 348.230 1073.590 349.410 1074.770 ;
        RECT 346.630 1071.990 347.810 1073.170 ;
        RECT 348.230 1071.990 349.410 1073.170 ;
        RECT 346.630 893.590 347.810 894.770 ;
        RECT 348.230 893.590 349.410 894.770 ;
        RECT 346.630 891.990 347.810 893.170 ;
        RECT 348.230 891.990 349.410 893.170 ;
        RECT 526.630 3558.160 527.810 3559.340 ;
        RECT 528.230 3558.160 529.410 3559.340 ;
        RECT 526.630 3556.560 527.810 3557.740 ;
        RECT 528.230 3556.560 529.410 3557.740 ;
        RECT 526.630 3413.590 527.810 3414.770 ;
        RECT 528.230 3413.590 529.410 3414.770 ;
        RECT 526.630 3411.990 527.810 3413.170 ;
        RECT 528.230 3411.990 529.410 3413.170 ;
        RECT 526.630 3233.590 527.810 3234.770 ;
        RECT 528.230 3233.590 529.410 3234.770 ;
        RECT 526.630 3231.990 527.810 3233.170 ;
        RECT 528.230 3231.990 529.410 3233.170 ;
        RECT 526.630 3053.590 527.810 3054.770 ;
        RECT 528.230 3053.590 529.410 3054.770 ;
        RECT 526.630 3051.990 527.810 3053.170 ;
        RECT 528.230 3051.990 529.410 3053.170 ;
        RECT 526.630 2873.590 527.810 2874.770 ;
        RECT 528.230 2873.590 529.410 2874.770 ;
        RECT 526.630 2871.990 527.810 2873.170 ;
        RECT 528.230 2871.990 529.410 2873.170 ;
        RECT 526.630 2693.590 527.810 2694.770 ;
        RECT 528.230 2693.590 529.410 2694.770 ;
        RECT 526.630 2691.990 527.810 2693.170 ;
        RECT 528.230 2691.990 529.410 2693.170 ;
        RECT 526.630 2513.590 527.810 2514.770 ;
        RECT 528.230 2513.590 529.410 2514.770 ;
        RECT 526.630 2511.990 527.810 2513.170 ;
        RECT 528.230 2511.990 529.410 2513.170 ;
        RECT 526.630 2333.590 527.810 2334.770 ;
        RECT 528.230 2333.590 529.410 2334.770 ;
        RECT 526.630 2331.990 527.810 2333.170 ;
        RECT 528.230 2331.990 529.410 2333.170 ;
        RECT 526.630 2153.590 527.810 2154.770 ;
        RECT 528.230 2153.590 529.410 2154.770 ;
        RECT 526.630 2151.990 527.810 2153.170 ;
        RECT 528.230 2151.990 529.410 2153.170 ;
        RECT 526.630 1973.590 527.810 1974.770 ;
        RECT 528.230 1973.590 529.410 1974.770 ;
        RECT 526.630 1971.990 527.810 1973.170 ;
        RECT 528.230 1971.990 529.410 1973.170 ;
        RECT 526.630 1793.590 527.810 1794.770 ;
        RECT 528.230 1793.590 529.410 1794.770 ;
        RECT 526.630 1791.990 527.810 1793.170 ;
        RECT 528.230 1791.990 529.410 1793.170 ;
        RECT 526.630 1613.590 527.810 1614.770 ;
        RECT 528.230 1613.590 529.410 1614.770 ;
        RECT 526.630 1611.990 527.810 1613.170 ;
        RECT 528.230 1611.990 529.410 1613.170 ;
        RECT 526.630 1433.590 527.810 1434.770 ;
        RECT 528.230 1433.590 529.410 1434.770 ;
        RECT 526.630 1431.990 527.810 1433.170 ;
        RECT 528.230 1431.990 529.410 1433.170 ;
        RECT 526.630 1253.590 527.810 1254.770 ;
        RECT 528.230 1253.590 529.410 1254.770 ;
        RECT 526.630 1251.990 527.810 1253.170 ;
        RECT 528.230 1251.990 529.410 1253.170 ;
        RECT 526.630 1073.590 527.810 1074.770 ;
        RECT 528.230 1073.590 529.410 1074.770 ;
        RECT 526.630 1071.990 527.810 1073.170 ;
        RECT 528.230 1071.990 529.410 1073.170 ;
        RECT 526.630 893.590 527.810 894.770 ;
        RECT 528.230 893.590 529.410 894.770 ;
        RECT 526.630 891.990 527.810 893.170 ;
        RECT 528.230 891.990 529.410 893.170 ;
        RECT 706.630 3558.160 707.810 3559.340 ;
        RECT 708.230 3558.160 709.410 3559.340 ;
        RECT 706.630 3556.560 707.810 3557.740 ;
        RECT 708.230 3556.560 709.410 3557.740 ;
        RECT 706.630 3413.590 707.810 3414.770 ;
        RECT 708.230 3413.590 709.410 3414.770 ;
        RECT 706.630 3411.990 707.810 3413.170 ;
        RECT 708.230 3411.990 709.410 3413.170 ;
        RECT 706.630 3233.590 707.810 3234.770 ;
        RECT 708.230 3233.590 709.410 3234.770 ;
        RECT 706.630 3231.990 707.810 3233.170 ;
        RECT 708.230 3231.990 709.410 3233.170 ;
        RECT 706.630 3053.590 707.810 3054.770 ;
        RECT 708.230 3053.590 709.410 3054.770 ;
        RECT 706.630 3051.990 707.810 3053.170 ;
        RECT 708.230 3051.990 709.410 3053.170 ;
        RECT 706.630 2873.590 707.810 2874.770 ;
        RECT 708.230 2873.590 709.410 2874.770 ;
        RECT 706.630 2871.990 707.810 2873.170 ;
        RECT 708.230 2871.990 709.410 2873.170 ;
        RECT 706.630 2693.590 707.810 2694.770 ;
        RECT 708.230 2693.590 709.410 2694.770 ;
        RECT 706.630 2691.990 707.810 2693.170 ;
        RECT 708.230 2691.990 709.410 2693.170 ;
        RECT 706.630 2513.590 707.810 2514.770 ;
        RECT 708.230 2513.590 709.410 2514.770 ;
        RECT 706.630 2511.990 707.810 2513.170 ;
        RECT 708.230 2511.990 709.410 2513.170 ;
        RECT 706.630 2333.590 707.810 2334.770 ;
        RECT 708.230 2333.590 709.410 2334.770 ;
        RECT 706.630 2331.990 707.810 2333.170 ;
        RECT 708.230 2331.990 709.410 2333.170 ;
        RECT 706.630 2153.590 707.810 2154.770 ;
        RECT 708.230 2153.590 709.410 2154.770 ;
        RECT 706.630 2151.990 707.810 2153.170 ;
        RECT 708.230 2151.990 709.410 2153.170 ;
        RECT 706.630 1973.590 707.810 1974.770 ;
        RECT 708.230 1973.590 709.410 1974.770 ;
        RECT 706.630 1971.990 707.810 1973.170 ;
        RECT 708.230 1971.990 709.410 1973.170 ;
        RECT 706.630 1793.590 707.810 1794.770 ;
        RECT 708.230 1793.590 709.410 1794.770 ;
        RECT 706.630 1791.990 707.810 1793.170 ;
        RECT 708.230 1791.990 709.410 1793.170 ;
        RECT 706.630 1613.590 707.810 1614.770 ;
        RECT 708.230 1613.590 709.410 1614.770 ;
        RECT 706.630 1611.990 707.810 1613.170 ;
        RECT 708.230 1611.990 709.410 1613.170 ;
        RECT 706.630 1433.590 707.810 1434.770 ;
        RECT 708.230 1433.590 709.410 1434.770 ;
        RECT 706.630 1431.990 707.810 1433.170 ;
        RECT 708.230 1431.990 709.410 1433.170 ;
        RECT 706.630 1253.590 707.810 1254.770 ;
        RECT 708.230 1253.590 709.410 1254.770 ;
        RECT 706.630 1251.990 707.810 1253.170 ;
        RECT 708.230 1251.990 709.410 1253.170 ;
        RECT 706.630 1073.590 707.810 1074.770 ;
        RECT 708.230 1073.590 709.410 1074.770 ;
        RECT 706.630 1071.990 707.810 1073.170 ;
        RECT 708.230 1071.990 709.410 1073.170 ;
        RECT 706.630 893.590 707.810 894.770 ;
        RECT 708.230 893.590 709.410 894.770 ;
        RECT 706.630 891.990 707.810 893.170 ;
        RECT 708.230 891.990 709.410 893.170 ;
        RECT 346.630 713.590 347.810 714.770 ;
        RECT 348.230 713.590 349.410 714.770 ;
        RECT 346.630 711.990 347.810 713.170 ;
        RECT 348.230 711.990 349.410 713.170 ;
        RECT 346.630 533.590 347.810 534.770 ;
        RECT 348.230 533.590 349.410 534.770 ;
        RECT 346.630 531.990 347.810 533.170 ;
        RECT 348.230 531.990 349.410 533.170 ;
        RECT 706.630 713.590 707.810 714.770 ;
        RECT 708.230 713.590 709.410 714.770 ;
        RECT 706.630 711.990 707.810 713.170 ;
        RECT 708.230 711.990 709.410 713.170 ;
        RECT 706.630 533.590 707.810 534.770 ;
        RECT 708.230 533.590 709.410 534.770 ;
        RECT 706.630 531.990 707.810 533.170 ;
        RECT 708.230 531.990 709.410 533.170 ;
        RECT 346.630 353.590 347.810 354.770 ;
        RECT 348.230 353.590 349.410 354.770 ;
        RECT 346.630 351.990 347.810 353.170 ;
        RECT 348.230 351.990 349.410 353.170 ;
        RECT 346.630 173.590 347.810 174.770 ;
        RECT 348.230 173.590 349.410 174.770 ;
        RECT 346.630 171.990 347.810 173.170 ;
        RECT 348.230 171.990 349.410 173.170 ;
        RECT 346.630 -38.060 347.810 -36.880 ;
        RECT 348.230 -38.060 349.410 -36.880 ;
        RECT 346.630 -39.660 347.810 -38.480 ;
        RECT 348.230 -39.660 349.410 -38.480 ;
        RECT 526.630 353.590 527.810 354.770 ;
        RECT 528.230 353.590 529.410 354.770 ;
        RECT 526.630 351.990 527.810 353.170 ;
        RECT 528.230 351.990 529.410 353.170 ;
        RECT 526.630 173.590 527.810 174.770 ;
        RECT 528.230 173.590 529.410 174.770 ;
        RECT 526.630 171.990 527.810 173.170 ;
        RECT 528.230 171.990 529.410 173.170 ;
        RECT 526.630 -38.060 527.810 -36.880 ;
        RECT 528.230 -38.060 529.410 -36.880 ;
        RECT 526.630 -39.660 527.810 -38.480 ;
        RECT 528.230 -39.660 529.410 -38.480 ;
        RECT 706.630 353.590 707.810 354.770 ;
        RECT 708.230 353.590 709.410 354.770 ;
        RECT 706.630 351.990 707.810 353.170 ;
        RECT 708.230 351.990 709.410 353.170 ;
        RECT 706.630 173.590 707.810 174.770 ;
        RECT 708.230 173.590 709.410 174.770 ;
        RECT 706.630 171.990 707.810 173.170 ;
        RECT 708.230 171.990 709.410 173.170 ;
        RECT 706.630 -38.060 707.810 -36.880 ;
        RECT 708.230 -38.060 709.410 -36.880 ;
        RECT 706.630 -39.660 707.810 -38.480 ;
        RECT 708.230 -39.660 709.410 -38.480 ;
        RECT 886.630 3558.160 887.810 3559.340 ;
        RECT 888.230 3558.160 889.410 3559.340 ;
        RECT 886.630 3556.560 887.810 3557.740 ;
        RECT 888.230 3556.560 889.410 3557.740 ;
        RECT 886.630 3413.590 887.810 3414.770 ;
        RECT 888.230 3413.590 889.410 3414.770 ;
        RECT 886.630 3411.990 887.810 3413.170 ;
        RECT 888.230 3411.990 889.410 3413.170 ;
        RECT 886.630 3233.590 887.810 3234.770 ;
        RECT 888.230 3233.590 889.410 3234.770 ;
        RECT 886.630 3231.990 887.810 3233.170 ;
        RECT 888.230 3231.990 889.410 3233.170 ;
        RECT 886.630 3053.590 887.810 3054.770 ;
        RECT 888.230 3053.590 889.410 3054.770 ;
        RECT 886.630 3051.990 887.810 3053.170 ;
        RECT 888.230 3051.990 889.410 3053.170 ;
        RECT 886.630 2873.590 887.810 2874.770 ;
        RECT 888.230 2873.590 889.410 2874.770 ;
        RECT 886.630 2871.990 887.810 2873.170 ;
        RECT 888.230 2871.990 889.410 2873.170 ;
        RECT 886.630 2693.590 887.810 2694.770 ;
        RECT 888.230 2693.590 889.410 2694.770 ;
        RECT 886.630 2691.990 887.810 2693.170 ;
        RECT 888.230 2691.990 889.410 2693.170 ;
        RECT 886.630 2513.590 887.810 2514.770 ;
        RECT 888.230 2513.590 889.410 2514.770 ;
        RECT 886.630 2511.990 887.810 2513.170 ;
        RECT 888.230 2511.990 889.410 2513.170 ;
        RECT 886.630 2333.590 887.810 2334.770 ;
        RECT 888.230 2333.590 889.410 2334.770 ;
        RECT 886.630 2331.990 887.810 2333.170 ;
        RECT 888.230 2331.990 889.410 2333.170 ;
        RECT 886.630 2153.590 887.810 2154.770 ;
        RECT 888.230 2153.590 889.410 2154.770 ;
        RECT 886.630 2151.990 887.810 2153.170 ;
        RECT 888.230 2151.990 889.410 2153.170 ;
        RECT 886.630 1973.590 887.810 1974.770 ;
        RECT 888.230 1973.590 889.410 1974.770 ;
        RECT 886.630 1971.990 887.810 1973.170 ;
        RECT 888.230 1971.990 889.410 1973.170 ;
        RECT 886.630 1793.590 887.810 1794.770 ;
        RECT 888.230 1793.590 889.410 1794.770 ;
        RECT 886.630 1791.990 887.810 1793.170 ;
        RECT 888.230 1791.990 889.410 1793.170 ;
        RECT 886.630 1613.590 887.810 1614.770 ;
        RECT 888.230 1613.590 889.410 1614.770 ;
        RECT 886.630 1611.990 887.810 1613.170 ;
        RECT 888.230 1611.990 889.410 1613.170 ;
        RECT 886.630 1433.590 887.810 1434.770 ;
        RECT 888.230 1433.590 889.410 1434.770 ;
        RECT 886.630 1431.990 887.810 1433.170 ;
        RECT 888.230 1431.990 889.410 1433.170 ;
        RECT 886.630 1253.590 887.810 1254.770 ;
        RECT 888.230 1253.590 889.410 1254.770 ;
        RECT 886.630 1251.990 887.810 1253.170 ;
        RECT 888.230 1251.990 889.410 1253.170 ;
        RECT 886.630 1073.590 887.810 1074.770 ;
        RECT 888.230 1073.590 889.410 1074.770 ;
        RECT 886.630 1071.990 887.810 1073.170 ;
        RECT 888.230 1071.990 889.410 1073.170 ;
        RECT 886.630 893.590 887.810 894.770 ;
        RECT 888.230 893.590 889.410 894.770 ;
        RECT 886.630 891.990 887.810 893.170 ;
        RECT 888.230 891.990 889.410 893.170 ;
        RECT 886.630 713.590 887.810 714.770 ;
        RECT 888.230 713.590 889.410 714.770 ;
        RECT 886.630 711.990 887.810 713.170 ;
        RECT 888.230 711.990 889.410 713.170 ;
        RECT 886.630 533.590 887.810 534.770 ;
        RECT 888.230 533.590 889.410 534.770 ;
        RECT 886.630 531.990 887.810 533.170 ;
        RECT 888.230 531.990 889.410 533.170 ;
        RECT 886.630 353.590 887.810 354.770 ;
        RECT 888.230 353.590 889.410 354.770 ;
        RECT 886.630 351.990 887.810 353.170 ;
        RECT 888.230 351.990 889.410 353.170 ;
        RECT 886.630 173.590 887.810 174.770 ;
        RECT 888.230 173.590 889.410 174.770 ;
        RECT 886.630 171.990 887.810 173.170 ;
        RECT 888.230 171.990 889.410 173.170 ;
        RECT 886.630 -38.060 887.810 -36.880 ;
        RECT 888.230 -38.060 889.410 -36.880 ;
        RECT 886.630 -39.660 887.810 -38.480 ;
        RECT 888.230 -39.660 889.410 -38.480 ;
        RECT 1066.630 3558.160 1067.810 3559.340 ;
        RECT 1068.230 3558.160 1069.410 3559.340 ;
        RECT 1066.630 3556.560 1067.810 3557.740 ;
        RECT 1068.230 3556.560 1069.410 3557.740 ;
        RECT 1066.630 3413.590 1067.810 3414.770 ;
        RECT 1068.230 3413.590 1069.410 3414.770 ;
        RECT 1066.630 3411.990 1067.810 3413.170 ;
        RECT 1068.230 3411.990 1069.410 3413.170 ;
        RECT 1066.630 3233.590 1067.810 3234.770 ;
        RECT 1068.230 3233.590 1069.410 3234.770 ;
        RECT 1066.630 3231.990 1067.810 3233.170 ;
        RECT 1068.230 3231.990 1069.410 3233.170 ;
        RECT 1066.630 3053.590 1067.810 3054.770 ;
        RECT 1068.230 3053.590 1069.410 3054.770 ;
        RECT 1066.630 3051.990 1067.810 3053.170 ;
        RECT 1068.230 3051.990 1069.410 3053.170 ;
        RECT 1066.630 2873.590 1067.810 2874.770 ;
        RECT 1068.230 2873.590 1069.410 2874.770 ;
        RECT 1066.630 2871.990 1067.810 2873.170 ;
        RECT 1068.230 2871.990 1069.410 2873.170 ;
        RECT 1066.630 2693.590 1067.810 2694.770 ;
        RECT 1068.230 2693.590 1069.410 2694.770 ;
        RECT 1066.630 2691.990 1067.810 2693.170 ;
        RECT 1068.230 2691.990 1069.410 2693.170 ;
        RECT 1066.630 2513.590 1067.810 2514.770 ;
        RECT 1068.230 2513.590 1069.410 2514.770 ;
        RECT 1066.630 2511.990 1067.810 2513.170 ;
        RECT 1068.230 2511.990 1069.410 2513.170 ;
        RECT 1066.630 2333.590 1067.810 2334.770 ;
        RECT 1068.230 2333.590 1069.410 2334.770 ;
        RECT 1066.630 2331.990 1067.810 2333.170 ;
        RECT 1068.230 2331.990 1069.410 2333.170 ;
        RECT 1066.630 2153.590 1067.810 2154.770 ;
        RECT 1068.230 2153.590 1069.410 2154.770 ;
        RECT 1066.630 2151.990 1067.810 2153.170 ;
        RECT 1068.230 2151.990 1069.410 2153.170 ;
        RECT 1066.630 1973.590 1067.810 1974.770 ;
        RECT 1068.230 1973.590 1069.410 1974.770 ;
        RECT 1066.630 1971.990 1067.810 1973.170 ;
        RECT 1068.230 1971.990 1069.410 1973.170 ;
        RECT 1066.630 1793.590 1067.810 1794.770 ;
        RECT 1068.230 1793.590 1069.410 1794.770 ;
        RECT 1066.630 1791.990 1067.810 1793.170 ;
        RECT 1068.230 1791.990 1069.410 1793.170 ;
        RECT 1066.630 1613.590 1067.810 1614.770 ;
        RECT 1068.230 1613.590 1069.410 1614.770 ;
        RECT 1066.630 1611.990 1067.810 1613.170 ;
        RECT 1068.230 1611.990 1069.410 1613.170 ;
        RECT 1066.630 1433.590 1067.810 1434.770 ;
        RECT 1068.230 1433.590 1069.410 1434.770 ;
        RECT 1066.630 1431.990 1067.810 1433.170 ;
        RECT 1068.230 1431.990 1069.410 1433.170 ;
        RECT 1066.630 1253.590 1067.810 1254.770 ;
        RECT 1068.230 1253.590 1069.410 1254.770 ;
        RECT 1066.630 1251.990 1067.810 1253.170 ;
        RECT 1068.230 1251.990 1069.410 1253.170 ;
        RECT 1066.630 1073.590 1067.810 1074.770 ;
        RECT 1068.230 1073.590 1069.410 1074.770 ;
        RECT 1066.630 1071.990 1067.810 1073.170 ;
        RECT 1068.230 1071.990 1069.410 1073.170 ;
        RECT 1066.630 893.590 1067.810 894.770 ;
        RECT 1068.230 893.590 1069.410 894.770 ;
        RECT 1066.630 891.990 1067.810 893.170 ;
        RECT 1068.230 891.990 1069.410 893.170 ;
        RECT 1066.630 713.590 1067.810 714.770 ;
        RECT 1068.230 713.590 1069.410 714.770 ;
        RECT 1066.630 711.990 1067.810 713.170 ;
        RECT 1068.230 711.990 1069.410 713.170 ;
        RECT 1066.630 533.590 1067.810 534.770 ;
        RECT 1068.230 533.590 1069.410 534.770 ;
        RECT 1066.630 531.990 1067.810 533.170 ;
        RECT 1068.230 531.990 1069.410 533.170 ;
        RECT 1066.630 353.590 1067.810 354.770 ;
        RECT 1068.230 353.590 1069.410 354.770 ;
        RECT 1066.630 351.990 1067.810 353.170 ;
        RECT 1068.230 351.990 1069.410 353.170 ;
        RECT 1066.630 173.590 1067.810 174.770 ;
        RECT 1068.230 173.590 1069.410 174.770 ;
        RECT 1066.630 171.990 1067.810 173.170 ;
        RECT 1068.230 171.990 1069.410 173.170 ;
        RECT 1066.630 -38.060 1067.810 -36.880 ;
        RECT 1068.230 -38.060 1069.410 -36.880 ;
        RECT 1066.630 -39.660 1067.810 -38.480 ;
        RECT 1068.230 -39.660 1069.410 -38.480 ;
        RECT 1246.630 3558.160 1247.810 3559.340 ;
        RECT 1248.230 3558.160 1249.410 3559.340 ;
        RECT 1246.630 3556.560 1247.810 3557.740 ;
        RECT 1248.230 3556.560 1249.410 3557.740 ;
        RECT 1246.630 3413.590 1247.810 3414.770 ;
        RECT 1248.230 3413.590 1249.410 3414.770 ;
        RECT 1246.630 3411.990 1247.810 3413.170 ;
        RECT 1248.230 3411.990 1249.410 3413.170 ;
        RECT 1246.630 3233.590 1247.810 3234.770 ;
        RECT 1248.230 3233.590 1249.410 3234.770 ;
        RECT 1246.630 3231.990 1247.810 3233.170 ;
        RECT 1248.230 3231.990 1249.410 3233.170 ;
        RECT 1246.630 3053.590 1247.810 3054.770 ;
        RECT 1248.230 3053.590 1249.410 3054.770 ;
        RECT 1246.630 3051.990 1247.810 3053.170 ;
        RECT 1248.230 3051.990 1249.410 3053.170 ;
        RECT 1246.630 2873.590 1247.810 2874.770 ;
        RECT 1248.230 2873.590 1249.410 2874.770 ;
        RECT 1246.630 2871.990 1247.810 2873.170 ;
        RECT 1248.230 2871.990 1249.410 2873.170 ;
        RECT 1246.630 2693.590 1247.810 2694.770 ;
        RECT 1248.230 2693.590 1249.410 2694.770 ;
        RECT 1246.630 2691.990 1247.810 2693.170 ;
        RECT 1248.230 2691.990 1249.410 2693.170 ;
        RECT 1246.630 2513.590 1247.810 2514.770 ;
        RECT 1248.230 2513.590 1249.410 2514.770 ;
        RECT 1246.630 2511.990 1247.810 2513.170 ;
        RECT 1248.230 2511.990 1249.410 2513.170 ;
        RECT 1246.630 2333.590 1247.810 2334.770 ;
        RECT 1248.230 2333.590 1249.410 2334.770 ;
        RECT 1246.630 2331.990 1247.810 2333.170 ;
        RECT 1248.230 2331.990 1249.410 2333.170 ;
        RECT 1246.630 2153.590 1247.810 2154.770 ;
        RECT 1248.230 2153.590 1249.410 2154.770 ;
        RECT 1246.630 2151.990 1247.810 2153.170 ;
        RECT 1248.230 2151.990 1249.410 2153.170 ;
        RECT 1246.630 1973.590 1247.810 1974.770 ;
        RECT 1248.230 1973.590 1249.410 1974.770 ;
        RECT 1246.630 1971.990 1247.810 1973.170 ;
        RECT 1248.230 1971.990 1249.410 1973.170 ;
        RECT 1246.630 1793.590 1247.810 1794.770 ;
        RECT 1248.230 1793.590 1249.410 1794.770 ;
        RECT 1246.630 1791.990 1247.810 1793.170 ;
        RECT 1248.230 1791.990 1249.410 1793.170 ;
        RECT 1246.630 1613.590 1247.810 1614.770 ;
        RECT 1248.230 1613.590 1249.410 1614.770 ;
        RECT 1246.630 1611.990 1247.810 1613.170 ;
        RECT 1248.230 1611.990 1249.410 1613.170 ;
        RECT 1246.630 1433.590 1247.810 1434.770 ;
        RECT 1248.230 1433.590 1249.410 1434.770 ;
        RECT 1246.630 1431.990 1247.810 1433.170 ;
        RECT 1248.230 1431.990 1249.410 1433.170 ;
        RECT 1246.630 1253.590 1247.810 1254.770 ;
        RECT 1248.230 1253.590 1249.410 1254.770 ;
        RECT 1246.630 1251.990 1247.810 1253.170 ;
        RECT 1248.230 1251.990 1249.410 1253.170 ;
        RECT 1246.630 1073.590 1247.810 1074.770 ;
        RECT 1248.230 1073.590 1249.410 1074.770 ;
        RECT 1246.630 1071.990 1247.810 1073.170 ;
        RECT 1248.230 1071.990 1249.410 1073.170 ;
        RECT 1246.630 893.590 1247.810 894.770 ;
        RECT 1248.230 893.590 1249.410 894.770 ;
        RECT 1246.630 891.990 1247.810 893.170 ;
        RECT 1248.230 891.990 1249.410 893.170 ;
        RECT 1246.630 713.590 1247.810 714.770 ;
        RECT 1248.230 713.590 1249.410 714.770 ;
        RECT 1246.630 711.990 1247.810 713.170 ;
        RECT 1248.230 711.990 1249.410 713.170 ;
        RECT 1246.630 533.590 1247.810 534.770 ;
        RECT 1248.230 533.590 1249.410 534.770 ;
        RECT 1246.630 531.990 1247.810 533.170 ;
        RECT 1248.230 531.990 1249.410 533.170 ;
        RECT 1246.630 353.590 1247.810 354.770 ;
        RECT 1248.230 353.590 1249.410 354.770 ;
        RECT 1246.630 351.990 1247.810 353.170 ;
        RECT 1248.230 351.990 1249.410 353.170 ;
        RECT 1246.630 173.590 1247.810 174.770 ;
        RECT 1248.230 173.590 1249.410 174.770 ;
        RECT 1246.630 171.990 1247.810 173.170 ;
        RECT 1248.230 171.990 1249.410 173.170 ;
        RECT 1246.630 -38.060 1247.810 -36.880 ;
        RECT 1248.230 -38.060 1249.410 -36.880 ;
        RECT 1246.630 -39.660 1247.810 -38.480 ;
        RECT 1248.230 -39.660 1249.410 -38.480 ;
        RECT 1426.630 3558.160 1427.810 3559.340 ;
        RECT 1428.230 3558.160 1429.410 3559.340 ;
        RECT 1426.630 3556.560 1427.810 3557.740 ;
        RECT 1428.230 3556.560 1429.410 3557.740 ;
        RECT 1426.630 3413.590 1427.810 3414.770 ;
        RECT 1428.230 3413.590 1429.410 3414.770 ;
        RECT 1426.630 3411.990 1427.810 3413.170 ;
        RECT 1428.230 3411.990 1429.410 3413.170 ;
        RECT 1426.630 3233.590 1427.810 3234.770 ;
        RECT 1428.230 3233.590 1429.410 3234.770 ;
        RECT 1426.630 3231.990 1427.810 3233.170 ;
        RECT 1428.230 3231.990 1429.410 3233.170 ;
        RECT 1426.630 3053.590 1427.810 3054.770 ;
        RECT 1428.230 3053.590 1429.410 3054.770 ;
        RECT 1426.630 3051.990 1427.810 3053.170 ;
        RECT 1428.230 3051.990 1429.410 3053.170 ;
        RECT 1426.630 2873.590 1427.810 2874.770 ;
        RECT 1428.230 2873.590 1429.410 2874.770 ;
        RECT 1426.630 2871.990 1427.810 2873.170 ;
        RECT 1428.230 2871.990 1429.410 2873.170 ;
        RECT 1426.630 2693.590 1427.810 2694.770 ;
        RECT 1428.230 2693.590 1429.410 2694.770 ;
        RECT 1426.630 2691.990 1427.810 2693.170 ;
        RECT 1428.230 2691.990 1429.410 2693.170 ;
        RECT 1426.630 2513.590 1427.810 2514.770 ;
        RECT 1428.230 2513.590 1429.410 2514.770 ;
        RECT 1426.630 2511.990 1427.810 2513.170 ;
        RECT 1428.230 2511.990 1429.410 2513.170 ;
        RECT 1426.630 2333.590 1427.810 2334.770 ;
        RECT 1428.230 2333.590 1429.410 2334.770 ;
        RECT 1426.630 2331.990 1427.810 2333.170 ;
        RECT 1428.230 2331.990 1429.410 2333.170 ;
        RECT 1426.630 2153.590 1427.810 2154.770 ;
        RECT 1428.230 2153.590 1429.410 2154.770 ;
        RECT 1426.630 2151.990 1427.810 2153.170 ;
        RECT 1428.230 2151.990 1429.410 2153.170 ;
        RECT 1426.630 1973.590 1427.810 1974.770 ;
        RECT 1428.230 1973.590 1429.410 1974.770 ;
        RECT 1426.630 1971.990 1427.810 1973.170 ;
        RECT 1428.230 1971.990 1429.410 1973.170 ;
        RECT 1426.630 1793.590 1427.810 1794.770 ;
        RECT 1428.230 1793.590 1429.410 1794.770 ;
        RECT 1426.630 1791.990 1427.810 1793.170 ;
        RECT 1428.230 1791.990 1429.410 1793.170 ;
        RECT 1426.630 1613.590 1427.810 1614.770 ;
        RECT 1428.230 1613.590 1429.410 1614.770 ;
        RECT 1426.630 1611.990 1427.810 1613.170 ;
        RECT 1428.230 1611.990 1429.410 1613.170 ;
        RECT 1426.630 1433.590 1427.810 1434.770 ;
        RECT 1428.230 1433.590 1429.410 1434.770 ;
        RECT 1426.630 1431.990 1427.810 1433.170 ;
        RECT 1428.230 1431.990 1429.410 1433.170 ;
        RECT 1426.630 1253.590 1427.810 1254.770 ;
        RECT 1428.230 1253.590 1429.410 1254.770 ;
        RECT 1426.630 1251.990 1427.810 1253.170 ;
        RECT 1428.230 1251.990 1429.410 1253.170 ;
        RECT 1426.630 1073.590 1427.810 1074.770 ;
        RECT 1428.230 1073.590 1429.410 1074.770 ;
        RECT 1426.630 1071.990 1427.810 1073.170 ;
        RECT 1428.230 1071.990 1429.410 1073.170 ;
        RECT 1426.630 893.590 1427.810 894.770 ;
        RECT 1428.230 893.590 1429.410 894.770 ;
        RECT 1426.630 891.990 1427.810 893.170 ;
        RECT 1428.230 891.990 1429.410 893.170 ;
        RECT 1426.630 713.590 1427.810 714.770 ;
        RECT 1428.230 713.590 1429.410 714.770 ;
        RECT 1426.630 711.990 1427.810 713.170 ;
        RECT 1428.230 711.990 1429.410 713.170 ;
        RECT 1426.630 533.590 1427.810 534.770 ;
        RECT 1428.230 533.590 1429.410 534.770 ;
        RECT 1426.630 531.990 1427.810 533.170 ;
        RECT 1428.230 531.990 1429.410 533.170 ;
        RECT 1426.630 353.590 1427.810 354.770 ;
        RECT 1428.230 353.590 1429.410 354.770 ;
        RECT 1426.630 351.990 1427.810 353.170 ;
        RECT 1428.230 351.990 1429.410 353.170 ;
        RECT 1426.630 173.590 1427.810 174.770 ;
        RECT 1428.230 173.590 1429.410 174.770 ;
        RECT 1426.630 171.990 1427.810 173.170 ;
        RECT 1428.230 171.990 1429.410 173.170 ;
        RECT 1426.630 -38.060 1427.810 -36.880 ;
        RECT 1428.230 -38.060 1429.410 -36.880 ;
        RECT 1426.630 -39.660 1427.810 -38.480 ;
        RECT 1428.230 -39.660 1429.410 -38.480 ;
        RECT 1606.630 3558.160 1607.810 3559.340 ;
        RECT 1608.230 3558.160 1609.410 3559.340 ;
        RECT 1606.630 3556.560 1607.810 3557.740 ;
        RECT 1608.230 3556.560 1609.410 3557.740 ;
        RECT 1606.630 3413.590 1607.810 3414.770 ;
        RECT 1608.230 3413.590 1609.410 3414.770 ;
        RECT 1606.630 3411.990 1607.810 3413.170 ;
        RECT 1608.230 3411.990 1609.410 3413.170 ;
        RECT 1606.630 3233.590 1607.810 3234.770 ;
        RECT 1608.230 3233.590 1609.410 3234.770 ;
        RECT 1606.630 3231.990 1607.810 3233.170 ;
        RECT 1608.230 3231.990 1609.410 3233.170 ;
        RECT 1606.630 3053.590 1607.810 3054.770 ;
        RECT 1608.230 3053.590 1609.410 3054.770 ;
        RECT 1606.630 3051.990 1607.810 3053.170 ;
        RECT 1608.230 3051.990 1609.410 3053.170 ;
        RECT 1606.630 2873.590 1607.810 2874.770 ;
        RECT 1608.230 2873.590 1609.410 2874.770 ;
        RECT 1606.630 2871.990 1607.810 2873.170 ;
        RECT 1608.230 2871.990 1609.410 2873.170 ;
        RECT 1606.630 2693.590 1607.810 2694.770 ;
        RECT 1608.230 2693.590 1609.410 2694.770 ;
        RECT 1606.630 2691.990 1607.810 2693.170 ;
        RECT 1608.230 2691.990 1609.410 2693.170 ;
        RECT 1606.630 2513.590 1607.810 2514.770 ;
        RECT 1608.230 2513.590 1609.410 2514.770 ;
        RECT 1606.630 2511.990 1607.810 2513.170 ;
        RECT 1608.230 2511.990 1609.410 2513.170 ;
        RECT 1606.630 2333.590 1607.810 2334.770 ;
        RECT 1608.230 2333.590 1609.410 2334.770 ;
        RECT 1606.630 2331.990 1607.810 2333.170 ;
        RECT 1608.230 2331.990 1609.410 2333.170 ;
        RECT 1606.630 2153.590 1607.810 2154.770 ;
        RECT 1608.230 2153.590 1609.410 2154.770 ;
        RECT 1606.630 2151.990 1607.810 2153.170 ;
        RECT 1608.230 2151.990 1609.410 2153.170 ;
        RECT 1606.630 1973.590 1607.810 1974.770 ;
        RECT 1608.230 1973.590 1609.410 1974.770 ;
        RECT 1606.630 1971.990 1607.810 1973.170 ;
        RECT 1608.230 1971.990 1609.410 1973.170 ;
        RECT 1606.630 1793.590 1607.810 1794.770 ;
        RECT 1608.230 1793.590 1609.410 1794.770 ;
        RECT 1606.630 1791.990 1607.810 1793.170 ;
        RECT 1608.230 1791.990 1609.410 1793.170 ;
        RECT 1606.630 1613.590 1607.810 1614.770 ;
        RECT 1608.230 1613.590 1609.410 1614.770 ;
        RECT 1606.630 1611.990 1607.810 1613.170 ;
        RECT 1608.230 1611.990 1609.410 1613.170 ;
        RECT 1606.630 1433.590 1607.810 1434.770 ;
        RECT 1608.230 1433.590 1609.410 1434.770 ;
        RECT 1606.630 1431.990 1607.810 1433.170 ;
        RECT 1608.230 1431.990 1609.410 1433.170 ;
        RECT 1606.630 1253.590 1607.810 1254.770 ;
        RECT 1608.230 1253.590 1609.410 1254.770 ;
        RECT 1606.630 1251.990 1607.810 1253.170 ;
        RECT 1608.230 1251.990 1609.410 1253.170 ;
        RECT 1606.630 1073.590 1607.810 1074.770 ;
        RECT 1608.230 1073.590 1609.410 1074.770 ;
        RECT 1606.630 1071.990 1607.810 1073.170 ;
        RECT 1608.230 1071.990 1609.410 1073.170 ;
        RECT 1606.630 893.590 1607.810 894.770 ;
        RECT 1608.230 893.590 1609.410 894.770 ;
        RECT 1606.630 891.990 1607.810 893.170 ;
        RECT 1608.230 891.990 1609.410 893.170 ;
        RECT 1606.630 713.590 1607.810 714.770 ;
        RECT 1608.230 713.590 1609.410 714.770 ;
        RECT 1606.630 711.990 1607.810 713.170 ;
        RECT 1608.230 711.990 1609.410 713.170 ;
        RECT 1606.630 533.590 1607.810 534.770 ;
        RECT 1608.230 533.590 1609.410 534.770 ;
        RECT 1606.630 531.990 1607.810 533.170 ;
        RECT 1608.230 531.990 1609.410 533.170 ;
        RECT 1606.630 353.590 1607.810 354.770 ;
        RECT 1608.230 353.590 1609.410 354.770 ;
        RECT 1606.630 351.990 1607.810 353.170 ;
        RECT 1608.230 351.990 1609.410 353.170 ;
        RECT 1606.630 173.590 1607.810 174.770 ;
        RECT 1608.230 173.590 1609.410 174.770 ;
        RECT 1606.630 171.990 1607.810 173.170 ;
        RECT 1608.230 171.990 1609.410 173.170 ;
        RECT 1606.630 -38.060 1607.810 -36.880 ;
        RECT 1608.230 -38.060 1609.410 -36.880 ;
        RECT 1606.630 -39.660 1607.810 -38.480 ;
        RECT 1608.230 -39.660 1609.410 -38.480 ;
        RECT 1786.630 3558.160 1787.810 3559.340 ;
        RECT 1788.230 3558.160 1789.410 3559.340 ;
        RECT 1786.630 3556.560 1787.810 3557.740 ;
        RECT 1788.230 3556.560 1789.410 3557.740 ;
        RECT 1786.630 3413.590 1787.810 3414.770 ;
        RECT 1788.230 3413.590 1789.410 3414.770 ;
        RECT 1786.630 3411.990 1787.810 3413.170 ;
        RECT 1788.230 3411.990 1789.410 3413.170 ;
        RECT 1786.630 3233.590 1787.810 3234.770 ;
        RECT 1788.230 3233.590 1789.410 3234.770 ;
        RECT 1786.630 3231.990 1787.810 3233.170 ;
        RECT 1788.230 3231.990 1789.410 3233.170 ;
        RECT 1786.630 3053.590 1787.810 3054.770 ;
        RECT 1788.230 3053.590 1789.410 3054.770 ;
        RECT 1786.630 3051.990 1787.810 3053.170 ;
        RECT 1788.230 3051.990 1789.410 3053.170 ;
        RECT 1786.630 2873.590 1787.810 2874.770 ;
        RECT 1788.230 2873.590 1789.410 2874.770 ;
        RECT 1786.630 2871.990 1787.810 2873.170 ;
        RECT 1788.230 2871.990 1789.410 2873.170 ;
        RECT 1786.630 2693.590 1787.810 2694.770 ;
        RECT 1788.230 2693.590 1789.410 2694.770 ;
        RECT 1786.630 2691.990 1787.810 2693.170 ;
        RECT 1788.230 2691.990 1789.410 2693.170 ;
        RECT 1786.630 2513.590 1787.810 2514.770 ;
        RECT 1788.230 2513.590 1789.410 2514.770 ;
        RECT 1786.630 2511.990 1787.810 2513.170 ;
        RECT 1788.230 2511.990 1789.410 2513.170 ;
        RECT 1786.630 2333.590 1787.810 2334.770 ;
        RECT 1788.230 2333.590 1789.410 2334.770 ;
        RECT 1786.630 2331.990 1787.810 2333.170 ;
        RECT 1788.230 2331.990 1789.410 2333.170 ;
        RECT 1786.630 2153.590 1787.810 2154.770 ;
        RECT 1788.230 2153.590 1789.410 2154.770 ;
        RECT 1786.630 2151.990 1787.810 2153.170 ;
        RECT 1788.230 2151.990 1789.410 2153.170 ;
        RECT 1786.630 1973.590 1787.810 1974.770 ;
        RECT 1788.230 1973.590 1789.410 1974.770 ;
        RECT 1786.630 1971.990 1787.810 1973.170 ;
        RECT 1788.230 1971.990 1789.410 1973.170 ;
        RECT 1786.630 1793.590 1787.810 1794.770 ;
        RECT 1788.230 1793.590 1789.410 1794.770 ;
        RECT 1786.630 1791.990 1787.810 1793.170 ;
        RECT 1788.230 1791.990 1789.410 1793.170 ;
        RECT 1786.630 1613.590 1787.810 1614.770 ;
        RECT 1788.230 1613.590 1789.410 1614.770 ;
        RECT 1786.630 1611.990 1787.810 1613.170 ;
        RECT 1788.230 1611.990 1789.410 1613.170 ;
        RECT 1786.630 1433.590 1787.810 1434.770 ;
        RECT 1788.230 1433.590 1789.410 1434.770 ;
        RECT 1786.630 1431.990 1787.810 1433.170 ;
        RECT 1788.230 1431.990 1789.410 1433.170 ;
        RECT 1786.630 1253.590 1787.810 1254.770 ;
        RECT 1788.230 1253.590 1789.410 1254.770 ;
        RECT 1786.630 1251.990 1787.810 1253.170 ;
        RECT 1788.230 1251.990 1789.410 1253.170 ;
        RECT 1786.630 1073.590 1787.810 1074.770 ;
        RECT 1788.230 1073.590 1789.410 1074.770 ;
        RECT 1786.630 1071.990 1787.810 1073.170 ;
        RECT 1788.230 1071.990 1789.410 1073.170 ;
        RECT 1786.630 893.590 1787.810 894.770 ;
        RECT 1788.230 893.590 1789.410 894.770 ;
        RECT 1786.630 891.990 1787.810 893.170 ;
        RECT 1788.230 891.990 1789.410 893.170 ;
        RECT 1786.630 713.590 1787.810 714.770 ;
        RECT 1788.230 713.590 1789.410 714.770 ;
        RECT 1786.630 711.990 1787.810 713.170 ;
        RECT 1788.230 711.990 1789.410 713.170 ;
        RECT 1786.630 533.590 1787.810 534.770 ;
        RECT 1788.230 533.590 1789.410 534.770 ;
        RECT 1786.630 531.990 1787.810 533.170 ;
        RECT 1788.230 531.990 1789.410 533.170 ;
        RECT 1786.630 353.590 1787.810 354.770 ;
        RECT 1788.230 353.590 1789.410 354.770 ;
        RECT 1786.630 351.990 1787.810 353.170 ;
        RECT 1788.230 351.990 1789.410 353.170 ;
        RECT 1786.630 173.590 1787.810 174.770 ;
        RECT 1788.230 173.590 1789.410 174.770 ;
        RECT 1786.630 171.990 1787.810 173.170 ;
        RECT 1788.230 171.990 1789.410 173.170 ;
        RECT 1786.630 -38.060 1787.810 -36.880 ;
        RECT 1788.230 -38.060 1789.410 -36.880 ;
        RECT 1786.630 -39.660 1787.810 -38.480 ;
        RECT 1788.230 -39.660 1789.410 -38.480 ;
        RECT 1966.630 3558.160 1967.810 3559.340 ;
        RECT 1968.230 3558.160 1969.410 3559.340 ;
        RECT 1966.630 3556.560 1967.810 3557.740 ;
        RECT 1968.230 3556.560 1969.410 3557.740 ;
        RECT 1966.630 3413.590 1967.810 3414.770 ;
        RECT 1968.230 3413.590 1969.410 3414.770 ;
        RECT 1966.630 3411.990 1967.810 3413.170 ;
        RECT 1968.230 3411.990 1969.410 3413.170 ;
        RECT 1966.630 3233.590 1967.810 3234.770 ;
        RECT 1968.230 3233.590 1969.410 3234.770 ;
        RECT 1966.630 3231.990 1967.810 3233.170 ;
        RECT 1968.230 3231.990 1969.410 3233.170 ;
        RECT 1966.630 3053.590 1967.810 3054.770 ;
        RECT 1968.230 3053.590 1969.410 3054.770 ;
        RECT 1966.630 3051.990 1967.810 3053.170 ;
        RECT 1968.230 3051.990 1969.410 3053.170 ;
        RECT 1966.630 2873.590 1967.810 2874.770 ;
        RECT 1968.230 2873.590 1969.410 2874.770 ;
        RECT 1966.630 2871.990 1967.810 2873.170 ;
        RECT 1968.230 2871.990 1969.410 2873.170 ;
        RECT 1966.630 2693.590 1967.810 2694.770 ;
        RECT 1968.230 2693.590 1969.410 2694.770 ;
        RECT 1966.630 2691.990 1967.810 2693.170 ;
        RECT 1968.230 2691.990 1969.410 2693.170 ;
        RECT 1966.630 2513.590 1967.810 2514.770 ;
        RECT 1968.230 2513.590 1969.410 2514.770 ;
        RECT 1966.630 2511.990 1967.810 2513.170 ;
        RECT 1968.230 2511.990 1969.410 2513.170 ;
        RECT 1966.630 2333.590 1967.810 2334.770 ;
        RECT 1968.230 2333.590 1969.410 2334.770 ;
        RECT 1966.630 2331.990 1967.810 2333.170 ;
        RECT 1968.230 2331.990 1969.410 2333.170 ;
        RECT 1966.630 2153.590 1967.810 2154.770 ;
        RECT 1968.230 2153.590 1969.410 2154.770 ;
        RECT 1966.630 2151.990 1967.810 2153.170 ;
        RECT 1968.230 2151.990 1969.410 2153.170 ;
        RECT 1966.630 1973.590 1967.810 1974.770 ;
        RECT 1968.230 1973.590 1969.410 1974.770 ;
        RECT 1966.630 1971.990 1967.810 1973.170 ;
        RECT 1968.230 1971.990 1969.410 1973.170 ;
        RECT 1966.630 1793.590 1967.810 1794.770 ;
        RECT 1968.230 1793.590 1969.410 1794.770 ;
        RECT 1966.630 1791.990 1967.810 1793.170 ;
        RECT 1968.230 1791.990 1969.410 1793.170 ;
        RECT 1966.630 1613.590 1967.810 1614.770 ;
        RECT 1968.230 1613.590 1969.410 1614.770 ;
        RECT 1966.630 1611.990 1967.810 1613.170 ;
        RECT 1968.230 1611.990 1969.410 1613.170 ;
        RECT 1966.630 1433.590 1967.810 1434.770 ;
        RECT 1968.230 1433.590 1969.410 1434.770 ;
        RECT 1966.630 1431.990 1967.810 1433.170 ;
        RECT 1968.230 1431.990 1969.410 1433.170 ;
        RECT 1966.630 1253.590 1967.810 1254.770 ;
        RECT 1968.230 1253.590 1969.410 1254.770 ;
        RECT 1966.630 1251.990 1967.810 1253.170 ;
        RECT 1968.230 1251.990 1969.410 1253.170 ;
        RECT 1966.630 1073.590 1967.810 1074.770 ;
        RECT 1968.230 1073.590 1969.410 1074.770 ;
        RECT 1966.630 1071.990 1967.810 1073.170 ;
        RECT 1968.230 1071.990 1969.410 1073.170 ;
        RECT 1966.630 893.590 1967.810 894.770 ;
        RECT 1968.230 893.590 1969.410 894.770 ;
        RECT 1966.630 891.990 1967.810 893.170 ;
        RECT 1968.230 891.990 1969.410 893.170 ;
        RECT 1966.630 713.590 1967.810 714.770 ;
        RECT 1968.230 713.590 1969.410 714.770 ;
        RECT 1966.630 711.990 1967.810 713.170 ;
        RECT 1968.230 711.990 1969.410 713.170 ;
        RECT 1966.630 533.590 1967.810 534.770 ;
        RECT 1968.230 533.590 1969.410 534.770 ;
        RECT 1966.630 531.990 1967.810 533.170 ;
        RECT 1968.230 531.990 1969.410 533.170 ;
        RECT 1966.630 353.590 1967.810 354.770 ;
        RECT 1968.230 353.590 1969.410 354.770 ;
        RECT 1966.630 351.990 1967.810 353.170 ;
        RECT 1968.230 351.990 1969.410 353.170 ;
        RECT 1966.630 173.590 1967.810 174.770 ;
        RECT 1968.230 173.590 1969.410 174.770 ;
        RECT 1966.630 171.990 1967.810 173.170 ;
        RECT 1968.230 171.990 1969.410 173.170 ;
        RECT 1966.630 -38.060 1967.810 -36.880 ;
        RECT 1968.230 -38.060 1969.410 -36.880 ;
        RECT 1966.630 -39.660 1967.810 -38.480 ;
        RECT 1968.230 -39.660 1969.410 -38.480 ;
        RECT 2146.630 3558.160 2147.810 3559.340 ;
        RECT 2148.230 3558.160 2149.410 3559.340 ;
        RECT 2146.630 3556.560 2147.810 3557.740 ;
        RECT 2148.230 3556.560 2149.410 3557.740 ;
        RECT 2146.630 3413.590 2147.810 3414.770 ;
        RECT 2148.230 3413.590 2149.410 3414.770 ;
        RECT 2146.630 3411.990 2147.810 3413.170 ;
        RECT 2148.230 3411.990 2149.410 3413.170 ;
        RECT 2146.630 3233.590 2147.810 3234.770 ;
        RECT 2148.230 3233.590 2149.410 3234.770 ;
        RECT 2146.630 3231.990 2147.810 3233.170 ;
        RECT 2148.230 3231.990 2149.410 3233.170 ;
        RECT 2146.630 3053.590 2147.810 3054.770 ;
        RECT 2148.230 3053.590 2149.410 3054.770 ;
        RECT 2146.630 3051.990 2147.810 3053.170 ;
        RECT 2148.230 3051.990 2149.410 3053.170 ;
        RECT 2146.630 2873.590 2147.810 2874.770 ;
        RECT 2148.230 2873.590 2149.410 2874.770 ;
        RECT 2146.630 2871.990 2147.810 2873.170 ;
        RECT 2148.230 2871.990 2149.410 2873.170 ;
        RECT 2146.630 2693.590 2147.810 2694.770 ;
        RECT 2148.230 2693.590 2149.410 2694.770 ;
        RECT 2146.630 2691.990 2147.810 2693.170 ;
        RECT 2148.230 2691.990 2149.410 2693.170 ;
        RECT 2146.630 2513.590 2147.810 2514.770 ;
        RECT 2148.230 2513.590 2149.410 2514.770 ;
        RECT 2146.630 2511.990 2147.810 2513.170 ;
        RECT 2148.230 2511.990 2149.410 2513.170 ;
        RECT 2146.630 2333.590 2147.810 2334.770 ;
        RECT 2148.230 2333.590 2149.410 2334.770 ;
        RECT 2146.630 2331.990 2147.810 2333.170 ;
        RECT 2148.230 2331.990 2149.410 2333.170 ;
        RECT 2146.630 2153.590 2147.810 2154.770 ;
        RECT 2148.230 2153.590 2149.410 2154.770 ;
        RECT 2146.630 2151.990 2147.810 2153.170 ;
        RECT 2148.230 2151.990 2149.410 2153.170 ;
        RECT 2146.630 1973.590 2147.810 1974.770 ;
        RECT 2148.230 1973.590 2149.410 1974.770 ;
        RECT 2146.630 1971.990 2147.810 1973.170 ;
        RECT 2148.230 1971.990 2149.410 1973.170 ;
        RECT 2146.630 1793.590 2147.810 1794.770 ;
        RECT 2148.230 1793.590 2149.410 1794.770 ;
        RECT 2146.630 1791.990 2147.810 1793.170 ;
        RECT 2148.230 1791.990 2149.410 1793.170 ;
        RECT 2146.630 1613.590 2147.810 1614.770 ;
        RECT 2148.230 1613.590 2149.410 1614.770 ;
        RECT 2146.630 1611.990 2147.810 1613.170 ;
        RECT 2148.230 1611.990 2149.410 1613.170 ;
        RECT 2146.630 1433.590 2147.810 1434.770 ;
        RECT 2148.230 1433.590 2149.410 1434.770 ;
        RECT 2146.630 1431.990 2147.810 1433.170 ;
        RECT 2148.230 1431.990 2149.410 1433.170 ;
        RECT 2146.630 1253.590 2147.810 1254.770 ;
        RECT 2148.230 1253.590 2149.410 1254.770 ;
        RECT 2146.630 1251.990 2147.810 1253.170 ;
        RECT 2148.230 1251.990 2149.410 1253.170 ;
        RECT 2146.630 1073.590 2147.810 1074.770 ;
        RECT 2148.230 1073.590 2149.410 1074.770 ;
        RECT 2146.630 1071.990 2147.810 1073.170 ;
        RECT 2148.230 1071.990 2149.410 1073.170 ;
        RECT 2146.630 893.590 2147.810 894.770 ;
        RECT 2148.230 893.590 2149.410 894.770 ;
        RECT 2146.630 891.990 2147.810 893.170 ;
        RECT 2148.230 891.990 2149.410 893.170 ;
        RECT 2146.630 713.590 2147.810 714.770 ;
        RECT 2148.230 713.590 2149.410 714.770 ;
        RECT 2146.630 711.990 2147.810 713.170 ;
        RECT 2148.230 711.990 2149.410 713.170 ;
        RECT 2146.630 533.590 2147.810 534.770 ;
        RECT 2148.230 533.590 2149.410 534.770 ;
        RECT 2146.630 531.990 2147.810 533.170 ;
        RECT 2148.230 531.990 2149.410 533.170 ;
        RECT 2146.630 353.590 2147.810 354.770 ;
        RECT 2148.230 353.590 2149.410 354.770 ;
        RECT 2146.630 351.990 2147.810 353.170 ;
        RECT 2148.230 351.990 2149.410 353.170 ;
        RECT 2146.630 173.590 2147.810 174.770 ;
        RECT 2148.230 173.590 2149.410 174.770 ;
        RECT 2146.630 171.990 2147.810 173.170 ;
        RECT 2148.230 171.990 2149.410 173.170 ;
        RECT 2146.630 -38.060 2147.810 -36.880 ;
        RECT 2148.230 -38.060 2149.410 -36.880 ;
        RECT 2146.630 -39.660 2147.810 -38.480 ;
        RECT 2148.230 -39.660 2149.410 -38.480 ;
        RECT 2326.630 3558.160 2327.810 3559.340 ;
        RECT 2328.230 3558.160 2329.410 3559.340 ;
        RECT 2326.630 3556.560 2327.810 3557.740 ;
        RECT 2328.230 3556.560 2329.410 3557.740 ;
        RECT 2326.630 3413.590 2327.810 3414.770 ;
        RECT 2328.230 3413.590 2329.410 3414.770 ;
        RECT 2326.630 3411.990 2327.810 3413.170 ;
        RECT 2328.230 3411.990 2329.410 3413.170 ;
        RECT 2326.630 3233.590 2327.810 3234.770 ;
        RECT 2328.230 3233.590 2329.410 3234.770 ;
        RECT 2326.630 3231.990 2327.810 3233.170 ;
        RECT 2328.230 3231.990 2329.410 3233.170 ;
        RECT 2326.630 3053.590 2327.810 3054.770 ;
        RECT 2328.230 3053.590 2329.410 3054.770 ;
        RECT 2326.630 3051.990 2327.810 3053.170 ;
        RECT 2328.230 3051.990 2329.410 3053.170 ;
        RECT 2326.630 2873.590 2327.810 2874.770 ;
        RECT 2328.230 2873.590 2329.410 2874.770 ;
        RECT 2326.630 2871.990 2327.810 2873.170 ;
        RECT 2328.230 2871.990 2329.410 2873.170 ;
        RECT 2326.630 2693.590 2327.810 2694.770 ;
        RECT 2328.230 2693.590 2329.410 2694.770 ;
        RECT 2326.630 2691.990 2327.810 2693.170 ;
        RECT 2328.230 2691.990 2329.410 2693.170 ;
        RECT 2326.630 2513.590 2327.810 2514.770 ;
        RECT 2328.230 2513.590 2329.410 2514.770 ;
        RECT 2326.630 2511.990 2327.810 2513.170 ;
        RECT 2328.230 2511.990 2329.410 2513.170 ;
        RECT 2326.630 2333.590 2327.810 2334.770 ;
        RECT 2328.230 2333.590 2329.410 2334.770 ;
        RECT 2326.630 2331.990 2327.810 2333.170 ;
        RECT 2328.230 2331.990 2329.410 2333.170 ;
        RECT 2326.630 2153.590 2327.810 2154.770 ;
        RECT 2328.230 2153.590 2329.410 2154.770 ;
        RECT 2326.630 2151.990 2327.810 2153.170 ;
        RECT 2328.230 2151.990 2329.410 2153.170 ;
        RECT 2326.630 1973.590 2327.810 1974.770 ;
        RECT 2328.230 1973.590 2329.410 1974.770 ;
        RECT 2326.630 1971.990 2327.810 1973.170 ;
        RECT 2328.230 1971.990 2329.410 1973.170 ;
        RECT 2326.630 1793.590 2327.810 1794.770 ;
        RECT 2328.230 1793.590 2329.410 1794.770 ;
        RECT 2326.630 1791.990 2327.810 1793.170 ;
        RECT 2328.230 1791.990 2329.410 1793.170 ;
        RECT 2326.630 1613.590 2327.810 1614.770 ;
        RECT 2328.230 1613.590 2329.410 1614.770 ;
        RECT 2326.630 1611.990 2327.810 1613.170 ;
        RECT 2328.230 1611.990 2329.410 1613.170 ;
        RECT 2326.630 1433.590 2327.810 1434.770 ;
        RECT 2328.230 1433.590 2329.410 1434.770 ;
        RECT 2326.630 1431.990 2327.810 1433.170 ;
        RECT 2328.230 1431.990 2329.410 1433.170 ;
        RECT 2326.630 1253.590 2327.810 1254.770 ;
        RECT 2328.230 1253.590 2329.410 1254.770 ;
        RECT 2326.630 1251.990 2327.810 1253.170 ;
        RECT 2328.230 1251.990 2329.410 1253.170 ;
        RECT 2326.630 1073.590 2327.810 1074.770 ;
        RECT 2328.230 1073.590 2329.410 1074.770 ;
        RECT 2326.630 1071.990 2327.810 1073.170 ;
        RECT 2328.230 1071.990 2329.410 1073.170 ;
        RECT 2326.630 893.590 2327.810 894.770 ;
        RECT 2328.230 893.590 2329.410 894.770 ;
        RECT 2326.630 891.990 2327.810 893.170 ;
        RECT 2328.230 891.990 2329.410 893.170 ;
        RECT 2326.630 713.590 2327.810 714.770 ;
        RECT 2328.230 713.590 2329.410 714.770 ;
        RECT 2326.630 711.990 2327.810 713.170 ;
        RECT 2328.230 711.990 2329.410 713.170 ;
        RECT 2326.630 533.590 2327.810 534.770 ;
        RECT 2328.230 533.590 2329.410 534.770 ;
        RECT 2326.630 531.990 2327.810 533.170 ;
        RECT 2328.230 531.990 2329.410 533.170 ;
        RECT 2326.630 353.590 2327.810 354.770 ;
        RECT 2328.230 353.590 2329.410 354.770 ;
        RECT 2326.630 351.990 2327.810 353.170 ;
        RECT 2328.230 351.990 2329.410 353.170 ;
        RECT 2326.630 173.590 2327.810 174.770 ;
        RECT 2328.230 173.590 2329.410 174.770 ;
        RECT 2326.630 171.990 2327.810 173.170 ;
        RECT 2328.230 171.990 2329.410 173.170 ;
        RECT 2326.630 -38.060 2327.810 -36.880 ;
        RECT 2328.230 -38.060 2329.410 -36.880 ;
        RECT 2326.630 -39.660 2327.810 -38.480 ;
        RECT 2328.230 -39.660 2329.410 -38.480 ;
        RECT 2506.630 3558.160 2507.810 3559.340 ;
        RECT 2508.230 3558.160 2509.410 3559.340 ;
        RECT 2506.630 3556.560 2507.810 3557.740 ;
        RECT 2508.230 3556.560 2509.410 3557.740 ;
        RECT 2506.630 3413.590 2507.810 3414.770 ;
        RECT 2508.230 3413.590 2509.410 3414.770 ;
        RECT 2506.630 3411.990 2507.810 3413.170 ;
        RECT 2508.230 3411.990 2509.410 3413.170 ;
        RECT 2506.630 3233.590 2507.810 3234.770 ;
        RECT 2508.230 3233.590 2509.410 3234.770 ;
        RECT 2506.630 3231.990 2507.810 3233.170 ;
        RECT 2508.230 3231.990 2509.410 3233.170 ;
        RECT 2506.630 3053.590 2507.810 3054.770 ;
        RECT 2508.230 3053.590 2509.410 3054.770 ;
        RECT 2506.630 3051.990 2507.810 3053.170 ;
        RECT 2508.230 3051.990 2509.410 3053.170 ;
        RECT 2506.630 2873.590 2507.810 2874.770 ;
        RECT 2508.230 2873.590 2509.410 2874.770 ;
        RECT 2506.630 2871.990 2507.810 2873.170 ;
        RECT 2508.230 2871.990 2509.410 2873.170 ;
        RECT 2506.630 2693.590 2507.810 2694.770 ;
        RECT 2508.230 2693.590 2509.410 2694.770 ;
        RECT 2506.630 2691.990 2507.810 2693.170 ;
        RECT 2508.230 2691.990 2509.410 2693.170 ;
        RECT 2506.630 2513.590 2507.810 2514.770 ;
        RECT 2508.230 2513.590 2509.410 2514.770 ;
        RECT 2506.630 2511.990 2507.810 2513.170 ;
        RECT 2508.230 2511.990 2509.410 2513.170 ;
        RECT 2506.630 2333.590 2507.810 2334.770 ;
        RECT 2508.230 2333.590 2509.410 2334.770 ;
        RECT 2506.630 2331.990 2507.810 2333.170 ;
        RECT 2508.230 2331.990 2509.410 2333.170 ;
        RECT 2506.630 2153.590 2507.810 2154.770 ;
        RECT 2508.230 2153.590 2509.410 2154.770 ;
        RECT 2506.630 2151.990 2507.810 2153.170 ;
        RECT 2508.230 2151.990 2509.410 2153.170 ;
        RECT 2506.630 1973.590 2507.810 1974.770 ;
        RECT 2508.230 1973.590 2509.410 1974.770 ;
        RECT 2506.630 1971.990 2507.810 1973.170 ;
        RECT 2508.230 1971.990 2509.410 1973.170 ;
        RECT 2506.630 1793.590 2507.810 1794.770 ;
        RECT 2508.230 1793.590 2509.410 1794.770 ;
        RECT 2506.630 1791.990 2507.810 1793.170 ;
        RECT 2508.230 1791.990 2509.410 1793.170 ;
        RECT 2506.630 1613.590 2507.810 1614.770 ;
        RECT 2508.230 1613.590 2509.410 1614.770 ;
        RECT 2506.630 1611.990 2507.810 1613.170 ;
        RECT 2508.230 1611.990 2509.410 1613.170 ;
        RECT 2506.630 1433.590 2507.810 1434.770 ;
        RECT 2508.230 1433.590 2509.410 1434.770 ;
        RECT 2506.630 1431.990 2507.810 1433.170 ;
        RECT 2508.230 1431.990 2509.410 1433.170 ;
        RECT 2506.630 1253.590 2507.810 1254.770 ;
        RECT 2508.230 1253.590 2509.410 1254.770 ;
        RECT 2506.630 1251.990 2507.810 1253.170 ;
        RECT 2508.230 1251.990 2509.410 1253.170 ;
        RECT 2506.630 1073.590 2507.810 1074.770 ;
        RECT 2508.230 1073.590 2509.410 1074.770 ;
        RECT 2506.630 1071.990 2507.810 1073.170 ;
        RECT 2508.230 1071.990 2509.410 1073.170 ;
        RECT 2506.630 893.590 2507.810 894.770 ;
        RECT 2508.230 893.590 2509.410 894.770 ;
        RECT 2506.630 891.990 2507.810 893.170 ;
        RECT 2508.230 891.990 2509.410 893.170 ;
        RECT 2506.630 713.590 2507.810 714.770 ;
        RECT 2508.230 713.590 2509.410 714.770 ;
        RECT 2506.630 711.990 2507.810 713.170 ;
        RECT 2508.230 711.990 2509.410 713.170 ;
        RECT 2506.630 533.590 2507.810 534.770 ;
        RECT 2508.230 533.590 2509.410 534.770 ;
        RECT 2506.630 531.990 2507.810 533.170 ;
        RECT 2508.230 531.990 2509.410 533.170 ;
        RECT 2506.630 353.590 2507.810 354.770 ;
        RECT 2508.230 353.590 2509.410 354.770 ;
        RECT 2506.630 351.990 2507.810 353.170 ;
        RECT 2508.230 351.990 2509.410 353.170 ;
        RECT 2506.630 173.590 2507.810 174.770 ;
        RECT 2508.230 173.590 2509.410 174.770 ;
        RECT 2506.630 171.990 2507.810 173.170 ;
        RECT 2508.230 171.990 2509.410 173.170 ;
        RECT 2506.630 -38.060 2507.810 -36.880 ;
        RECT 2508.230 -38.060 2509.410 -36.880 ;
        RECT 2506.630 -39.660 2507.810 -38.480 ;
        RECT 2508.230 -39.660 2509.410 -38.480 ;
        RECT 2686.630 3558.160 2687.810 3559.340 ;
        RECT 2688.230 3558.160 2689.410 3559.340 ;
        RECT 2686.630 3556.560 2687.810 3557.740 ;
        RECT 2688.230 3556.560 2689.410 3557.740 ;
        RECT 2686.630 3413.590 2687.810 3414.770 ;
        RECT 2688.230 3413.590 2689.410 3414.770 ;
        RECT 2686.630 3411.990 2687.810 3413.170 ;
        RECT 2688.230 3411.990 2689.410 3413.170 ;
        RECT 2686.630 3233.590 2687.810 3234.770 ;
        RECT 2688.230 3233.590 2689.410 3234.770 ;
        RECT 2686.630 3231.990 2687.810 3233.170 ;
        RECT 2688.230 3231.990 2689.410 3233.170 ;
        RECT 2686.630 3053.590 2687.810 3054.770 ;
        RECT 2688.230 3053.590 2689.410 3054.770 ;
        RECT 2686.630 3051.990 2687.810 3053.170 ;
        RECT 2688.230 3051.990 2689.410 3053.170 ;
        RECT 2686.630 2873.590 2687.810 2874.770 ;
        RECT 2688.230 2873.590 2689.410 2874.770 ;
        RECT 2686.630 2871.990 2687.810 2873.170 ;
        RECT 2688.230 2871.990 2689.410 2873.170 ;
        RECT 2686.630 2693.590 2687.810 2694.770 ;
        RECT 2688.230 2693.590 2689.410 2694.770 ;
        RECT 2686.630 2691.990 2687.810 2693.170 ;
        RECT 2688.230 2691.990 2689.410 2693.170 ;
        RECT 2686.630 2513.590 2687.810 2514.770 ;
        RECT 2688.230 2513.590 2689.410 2514.770 ;
        RECT 2686.630 2511.990 2687.810 2513.170 ;
        RECT 2688.230 2511.990 2689.410 2513.170 ;
        RECT 2686.630 2333.590 2687.810 2334.770 ;
        RECT 2688.230 2333.590 2689.410 2334.770 ;
        RECT 2686.630 2331.990 2687.810 2333.170 ;
        RECT 2688.230 2331.990 2689.410 2333.170 ;
        RECT 2686.630 2153.590 2687.810 2154.770 ;
        RECT 2688.230 2153.590 2689.410 2154.770 ;
        RECT 2686.630 2151.990 2687.810 2153.170 ;
        RECT 2688.230 2151.990 2689.410 2153.170 ;
        RECT 2686.630 1973.590 2687.810 1974.770 ;
        RECT 2688.230 1973.590 2689.410 1974.770 ;
        RECT 2686.630 1971.990 2687.810 1973.170 ;
        RECT 2688.230 1971.990 2689.410 1973.170 ;
        RECT 2686.630 1793.590 2687.810 1794.770 ;
        RECT 2688.230 1793.590 2689.410 1794.770 ;
        RECT 2686.630 1791.990 2687.810 1793.170 ;
        RECT 2688.230 1791.990 2689.410 1793.170 ;
        RECT 2686.630 1613.590 2687.810 1614.770 ;
        RECT 2688.230 1613.590 2689.410 1614.770 ;
        RECT 2686.630 1611.990 2687.810 1613.170 ;
        RECT 2688.230 1611.990 2689.410 1613.170 ;
        RECT 2686.630 1433.590 2687.810 1434.770 ;
        RECT 2688.230 1433.590 2689.410 1434.770 ;
        RECT 2686.630 1431.990 2687.810 1433.170 ;
        RECT 2688.230 1431.990 2689.410 1433.170 ;
        RECT 2686.630 1253.590 2687.810 1254.770 ;
        RECT 2688.230 1253.590 2689.410 1254.770 ;
        RECT 2686.630 1251.990 2687.810 1253.170 ;
        RECT 2688.230 1251.990 2689.410 1253.170 ;
        RECT 2686.630 1073.590 2687.810 1074.770 ;
        RECT 2688.230 1073.590 2689.410 1074.770 ;
        RECT 2686.630 1071.990 2687.810 1073.170 ;
        RECT 2688.230 1071.990 2689.410 1073.170 ;
        RECT 2686.630 893.590 2687.810 894.770 ;
        RECT 2688.230 893.590 2689.410 894.770 ;
        RECT 2686.630 891.990 2687.810 893.170 ;
        RECT 2688.230 891.990 2689.410 893.170 ;
        RECT 2686.630 713.590 2687.810 714.770 ;
        RECT 2688.230 713.590 2689.410 714.770 ;
        RECT 2686.630 711.990 2687.810 713.170 ;
        RECT 2688.230 711.990 2689.410 713.170 ;
        RECT 2686.630 533.590 2687.810 534.770 ;
        RECT 2688.230 533.590 2689.410 534.770 ;
        RECT 2686.630 531.990 2687.810 533.170 ;
        RECT 2688.230 531.990 2689.410 533.170 ;
        RECT 2686.630 353.590 2687.810 354.770 ;
        RECT 2688.230 353.590 2689.410 354.770 ;
        RECT 2686.630 351.990 2687.810 353.170 ;
        RECT 2688.230 351.990 2689.410 353.170 ;
        RECT 2686.630 173.590 2687.810 174.770 ;
        RECT 2688.230 173.590 2689.410 174.770 ;
        RECT 2686.630 171.990 2687.810 173.170 ;
        RECT 2688.230 171.990 2689.410 173.170 ;
        RECT 2686.630 -38.060 2687.810 -36.880 ;
        RECT 2688.230 -38.060 2689.410 -36.880 ;
        RECT 2686.630 -39.660 2687.810 -38.480 ;
        RECT 2688.230 -39.660 2689.410 -38.480 ;
        RECT 2866.630 3558.160 2867.810 3559.340 ;
        RECT 2868.230 3558.160 2869.410 3559.340 ;
        RECT 2866.630 3556.560 2867.810 3557.740 ;
        RECT 2868.230 3556.560 2869.410 3557.740 ;
        RECT 2866.630 3413.590 2867.810 3414.770 ;
        RECT 2868.230 3413.590 2869.410 3414.770 ;
        RECT 2866.630 3411.990 2867.810 3413.170 ;
        RECT 2868.230 3411.990 2869.410 3413.170 ;
        RECT 2866.630 3233.590 2867.810 3234.770 ;
        RECT 2868.230 3233.590 2869.410 3234.770 ;
        RECT 2866.630 3231.990 2867.810 3233.170 ;
        RECT 2868.230 3231.990 2869.410 3233.170 ;
        RECT 2866.630 3053.590 2867.810 3054.770 ;
        RECT 2868.230 3053.590 2869.410 3054.770 ;
        RECT 2866.630 3051.990 2867.810 3053.170 ;
        RECT 2868.230 3051.990 2869.410 3053.170 ;
        RECT 2866.630 2873.590 2867.810 2874.770 ;
        RECT 2868.230 2873.590 2869.410 2874.770 ;
        RECT 2866.630 2871.990 2867.810 2873.170 ;
        RECT 2868.230 2871.990 2869.410 2873.170 ;
        RECT 2866.630 2693.590 2867.810 2694.770 ;
        RECT 2868.230 2693.590 2869.410 2694.770 ;
        RECT 2866.630 2691.990 2867.810 2693.170 ;
        RECT 2868.230 2691.990 2869.410 2693.170 ;
        RECT 2866.630 2513.590 2867.810 2514.770 ;
        RECT 2868.230 2513.590 2869.410 2514.770 ;
        RECT 2866.630 2511.990 2867.810 2513.170 ;
        RECT 2868.230 2511.990 2869.410 2513.170 ;
        RECT 2866.630 2333.590 2867.810 2334.770 ;
        RECT 2868.230 2333.590 2869.410 2334.770 ;
        RECT 2866.630 2331.990 2867.810 2333.170 ;
        RECT 2868.230 2331.990 2869.410 2333.170 ;
        RECT 2866.630 2153.590 2867.810 2154.770 ;
        RECT 2868.230 2153.590 2869.410 2154.770 ;
        RECT 2866.630 2151.990 2867.810 2153.170 ;
        RECT 2868.230 2151.990 2869.410 2153.170 ;
        RECT 2866.630 1973.590 2867.810 1974.770 ;
        RECT 2868.230 1973.590 2869.410 1974.770 ;
        RECT 2866.630 1971.990 2867.810 1973.170 ;
        RECT 2868.230 1971.990 2869.410 1973.170 ;
        RECT 2866.630 1793.590 2867.810 1794.770 ;
        RECT 2868.230 1793.590 2869.410 1794.770 ;
        RECT 2866.630 1791.990 2867.810 1793.170 ;
        RECT 2868.230 1791.990 2869.410 1793.170 ;
        RECT 2866.630 1613.590 2867.810 1614.770 ;
        RECT 2868.230 1613.590 2869.410 1614.770 ;
        RECT 2866.630 1611.990 2867.810 1613.170 ;
        RECT 2868.230 1611.990 2869.410 1613.170 ;
        RECT 2866.630 1433.590 2867.810 1434.770 ;
        RECT 2868.230 1433.590 2869.410 1434.770 ;
        RECT 2866.630 1431.990 2867.810 1433.170 ;
        RECT 2868.230 1431.990 2869.410 1433.170 ;
        RECT 2866.630 1253.590 2867.810 1254.770 ;
        RECT 2868.230 1253.590 2869.410 1254.770 ;
        RECT 2866.630 1251.990 2867.810 1253.170 ;
        RECT 2868.230 1251.990 2869.410 1253.170 ;
        RECT 2866.630 1073.590 2867.810 1074.770 ;
        RECT 2868.230 1073.590 2869.410 1074.770 ;
        RECT 2866.630 1071.990 2867.810 1073.170 ;
        RECT 2868.230 1071.990 2869.410 1073.170 ;
        RECT 2866.630 893.590 2867.810 894.770 ;
        RECT 2868.230 893.590 2869.410 894.770 ;
        RECT 2866.630 891.990 2867.810 893.170 ;
        RECT 2868.230 891.990 2869.410 893.170 ;
        RECT 2866.630 713.590 2867.810 714.770 ;
        RECT 2868.230 713.590 2869.410 714.770 ;
        RECT 2866.630 711.990 2867.810 713.170 ;
        RECT 2868.230 711.990 2869.410 713.170 ;
        RECT 2866.630 533.590 2867.810 534.770 ;
        RECT 2868.230 533.590 2869.410 534.770 ;
        RECT 2866.630 531.990 2867.810 533.170 ;
        RECT 2868.230 531.990 2869.410 533.170 ;
        RECT 2866.630 353.590 2867.810 354.770 ;
        RECT 2868.230 353.590 2869.410 354.770 ;
        RECT 2866.630 351.990 2867.810 353.170 ;
        RECT 2868.230 351.990 2869.410 353.170 ;
        RECT 2866.630 173.590 2867.810 174.770 ;
        RECT 2868.230 173.590 2869.410 174.770 ;
        RECT 2866.630 171.990 2867.810 173.170 ;
        RECT 2868.230 171.990 2869.410 173.170 ;
        RECT 2866.630 -38.060 2867.810 -36.880 ;
        RECT 2868.230 -38.060 2869.410 -36.880 ;
        RECT 2866.630 -39.660 2867.810 -38.480 ;
        RECT 2868.230 -39.660 2869.410 -38.480 ;
        RECT 2961.860 3558.160 2963.040 3559.340 ;
        RECT 2963.460 3558.160 2964.640 3559.340 ;
        RECT 2961.860 3556.560 2963.040 3557.740 ;
        RECT 2963.460 3556.560 2964.640 3557.740 ;
        RECT 2961.860 3413.590 2963.040 3414.770 ;
        RECT 2963.460 3413.590 2964.640 3414.770 ;
        RECT 2961.860 3411.990 2963.040 3413.170 ;
        RECT 2963.460 3411.990 2964.640 3413.170 ;
        RECT 2961.860 3233.590 2963.040 3234.770 ;
        RECT 2963.460 3233.590 2964.640 3234.770 ;
        RECT 2961.860 3231.990 2963.040 3233.170 ;
        RECT 2963.460 3231.990 2964.640 3233.170 ;
        RECT 2961.860 3053.590 2963.040 3054.770 ;
        RECT 2963.460 3053.590 2964.640 3054.770 ;
        RECT 2961.860 3051.990 2963.040 3053.170 ;
        RECT 2963.460 3051.990 2964.640 3053.170 ;
        RECT 2961.860 2873.590 2963.040 2874.770 ;
        RECT 2963.460 2873.590 2964.640 2874.770 ;
        RECT 2961.860 2871.990 2963.040 2873.170 ;
        RECT 2963.460 2871.990 2964.640 2873.170 ;
        RECT 2961.860 2693.590 2963.040 2694.770 ;
        RECT 2963.460 2693.590 2964.640 2694.770 ;
        RECT 2961.860 2691.990 2963.040 2693.170 ;
        RECT 2963.460 2691.990 2964.640 2693.170 ;
        RECT 2961.860 2513.590 2963.040 2514.770 ;
        RECT 2963.460 2513.590 2964.640 2514.770 ;
        RECT 2961.860 2511.990 2963.040 2513.170 ;
        RECT 2963.460 2511.990 2964.640 2513.170 ;
        RECT 2961.860 2333.590 2963.040 2334.770 ;
        RECT 2963.460 2333.590 2964.640 2334.770 ;
        RECT 2961.860 2331.990 2963.040 2333.170 ;
        RECT 2963.460 2331.990 2964.640 2333.170 ;
        RECT 2961.860 2153.590 2963.040 2154.770 ;
        RECT 2963.460 2153.590 2964.640 2154.770 ;
        RECT 2961.860 2151.990 2963.040 2153.170 ;
        RECT 2963.460 2151.990 2964.640 2153.170 ;
        RECT 2961.860 1973.590 2963.040 1974.770 ;
        RECT 2963.460 1973.590 2964.640 1974.770 ;
        RECT 2961.860 1971.990 2963.040 1973.170 ;
        RECT 2963.460 1971.990 2964.640 1973.170 ;
        RECT 2961.860 1793.590 2963.040 1794.770 ;
        RECT 2963.460 1793.590 2964.640 1794.770 ;
        RECT 2961.860 1791.990 2963.040 1793.170 ;
        RECT 2963.460 1791.990 2964.640 1793.170 ;
        RECT 2961.860 1613.590 2963.040 1614.770 ;
        RECT 2963.460 1613.590 2964.640 1614.770 ;
        RECT 2961.860 1611.990 2963.040 1613.170 ;
        RECT 2963.460 1611.990 2964.640 1613.170 ;
        RECT 2961.860 1433.590 2963.040 1434.770 ;
        RECT 2963.460 1433.590 2964.640 1434.770 ;
        RECT 2961.860 1431.990 2963.040 1433.170 ;
        RECT 2963.460 1431.990 2964.640 1433.170 ;
        RECT 2961.860 1253.590 2963.040 1254.770 ;
        RECT 2963.460 1253.590 2964.640 1254.770 ;
        RECT 2961.860 1251.990 2963.040 1253.170 ;
        RECT 2963.460 1251.990 2964.640 1253.170 ;
        RECT 2961.860 1073.590 2963.040 1074.770 ;
        RECT 2963.460 1073.590 2964.640 1074.770 ;
        RECT 2961.860 1071.990 2963.040 1073.170 ;
        RECT 2963.460 1071.990 2964.640 1073.170 ;
        RECT 2961.860 893.590 2963.040 894.770 ;
        RECT 2963.460 893.590 2964.640 894.770 ;
        RECT 2961.860 891.990 2963.040 893.170 ;
        RECT 2963.460 891.990 2964.640 893.170 ;
        RECT 2961.860 713.590 2963.040 714.770 ;
        RECT 2963.460 713.590 2964.640 714.770 ;
        RECT 2961.860 711.990 2963.040 713.170 ;
        RECT 2963.460 711.990 2964.640 713.170 ;
        RECT 2961.860 533.590 2963.040 534.770 ;
        RECT 2963.460 533.590 2964.640 534.770 ;
        RECT 2961.860 531.990 2963.040 533.170 ;
        RECT 2963.460 531.990 2964.640 533.170 ;
        RECT 2961.860 353.590 2963.040 354.770 ;
        RECT 2963.460 353.590 2964.640 354.770 ;
        RECT 2961.860 351.990 2963.040 353.170 ;
        RECT 2963.460 351.990 2964.640 353.170 ;
        RECT 2961.860 173.590 2963.040 174.770 ;
        RECT 2963.460 173.590 2964.640 174.770 ;
        RECT 2961.860 171.990 2963.040 173.170 ;
        RECT 2963.460 171.990 2964.640 173.170 ;
        RECT 2961.860 -38.060 2963.040 -36.880 ;
        RECT 2963.460 -38.060 2964.640 -36.880 ;
        RECT 2961.860 -39.660 2963.040 -38.480 ;
        RECT 2963.460 -39.660 2964.640 -38.480 ;
      LAYER met5 ;
        RECT -45.180 3556.400 2964.800 3559.500 ;
        RECT -45.180 3411.830 2964.800 3414.930 ;
        RECT -45.180 3231.830 2964.800 3234.930 ;
        RECT -45.180 3051.830 2964.800 3054.930 ;
        RECT -45.180 2871.830 2964.800 2874.930 ;
        RECT -45.180 2691.830 2964.800 2694.930 ;
        RECT -45.180 2511.830 2964.800 2514.930 ;
        RECT -45.180 2331.830 2964.800 2334.930 ;
        RECT -45.180 2151.830 2964.800 2154.930 ;
        RECT -45.180 1971.830 2964.800 1974.930 ;
        RECT -45.180 1791.830 2964.800 1794.930 ;
        RECT -45.180 1611.830 2964.800 1614.930 ;
        RECT -45.180 1431.830 2964.800 1434.930 ;
        RECT -45.180 1251.830 2964.800 1254.930 ;
        RECT -45.180 1071.830 2964.800 1074.930 ;
        RECT -45.180 891.830 2964.800 894.930 ;
        RECT -45.180 711.830 2964.800 714.930 ;
        RECT -45.180 531.830 2964.800 534.930 ;
        RECT -45.180 351.830 2964.800 354.930 ;
        RECT -45.180 171.830 2964.800 174.930 ;
        RECT -45.180 -39.820 2964.800 -36.720 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
        RECT 31.470 -39.820 34.570 3559.500 ;
        RECT 211.470 -39.820 214.570 3559.500 ;
        RECT 391.470 760.000 394.570 3559.500 ;
        RECT 571.470 760.000 574.570 3559.500 ;
        RECT 497.840 510.640 499.440 736.880 ;
        RECT 391.470 -39.820 394.570 490.000 ;
        RECT 571.470 -39.820 574.570 490.000 ;
        RECT 751.470 -39.820 754.570 3559.500 ;
        RECT 931.470 -39.820 934.570 3559.500 ;
        RECT 1111.470 -39.820 1114.570 3559.500 ;
        RECT 1291.470 -39.820 1294.570 3559.500 ;
        RECT 1471.470 -39.820 1474.570 3559.500 ;
        RECT 1651.470 -39.820 1654.570 3559.500 ;
        RECT 1831.470 -39.820 1834.570 3559.500 ;
        RECT 2011.470 -39.820 2014.570 3559.500 ;
        RECT 2191.470 -39.820 2194.570 3559.500 ;
        RECT 2371.470 -39.820 2374.570 3559.500 ;
        RECT 2551.470 -39.820 2554.570 3559.500 ;
        RECT 2731.470 -39.820 2734.570 3559.500 ;
        RECT 2911.470 -39.820 2914.570 3559.500 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
      LAYER via4 ;
        RECT -16.220 3529.360 -15.040 3530.540 ;
        RECT -14.620 3529.360 -13.440 3530.540 ;
        RECT -16.220 3527.760 -15.040 3528.940 ;
        RECT -14.620 3527.760 -13.440 3528.940 ;
        RECT -16.220 3458.590 -15.040 3459.770 ;
        RECT -14.620 3458.590 -13.440 3459.770 ;
        RECT -16.220 3456.990 -15.040 3458.170 ;
        RECT -14.620 3456.990 -13.440 3458.170 ;
        RECT -16.220 3278.590 -15.040 3279.770 ;
        RECT -14.620 3278.590 -13.440 3279.770 ;
        RECT -16.220 3276.990 -15.040 3278.170 ;
        RECT -14.620 3276.990 -13.440 3278.170 ;
        RECT -16.220 3098.590 -15.040 3099.770 ;
        RECT -14.620 3098.590 -13.440 3099.770 ;
        RECT -16.220 3096.990 -15.040 3098.170 ;
        RECT -14.620 3096.990 -13.440 3098.170 ;
        RECT -16.220 2918.590 -15.040 2919.770 ;
        RECT -14.620 2918.590 -13.440 2919.770 ;
        RECT -16.220 2916.990 -15.040 2918.170 ;
        RECT -14.620 2916.990 -13.440 2918.170 ;
        RECT -16.220 2738.590 -15.040 2739.770 ;
        RECT -14.620 2738.590 -13.440 2739.770 ;
        RECT -16.220 2736.990 -15.040 2738.170 ;
        RECT -14.620 2736.990 -13.440 2738.170 ;
        RECT -16.220 2558.590 -15.040 2559.770 ;
        RECT -14.620 2558.590 -13.440 2559.770 ;
        RECT -16.220 2556.990 -15.040 2558.170 ;
        RECT -14.620 2556.990 -13.440 2558.170 ;
        RECT -16.220 2378.590 -15.040 2379.770 ;
        RECT -14.620 2378.590 -13.440 2379.770 ;
        RECT -16.220 2376.990 -15.040 2378.170 ;
        RECT -14.620 2376.990 -13.440 2378.170 ;
        RECT -16.220 2198.590 -15.040 2199.770 ;
        RECT -14.620 2198.590 -13.440 2199.770 ;
        RECT -16.220 2196.990 -15.040 2198.170 ;
        RECT -14.620 2196.990 -13.440 2198.170 ;
        RECT -16.220 2018.590 -15.040 2019.770 ;
        RECT -14.620 2018.590 -13.440 2019.770 ;
        RECT -16.220 2016.990 -15.040 2018.170 ;
        RECT -14.620 2016.990 -13.440 2018.170 ;
        RECT -16.220 1838.590 -15.040 1839.770 ;
        RECT -14.620 1838.590 -13.440 1839.770 ;
        RECT -16.220 1836.990 -15.040 1838.170 ;
        RECT -14.620 1836.990 -13.440 1838.170 ;
        RECT -16.220 1658.590 -15.040 1659.770 ;
        RECT -14.620 1658.590 -13.440 1659.770 ;
        RECT -16.220 1656.990 -15.040 1658.170 ;
        RECT -14.620 1656.990 -13.440 1658.170 ;
        RECT -16.220 1478.590 -15.040 1479.770 ;
        RECT -14.620 1478.590 -13.440 1479.770 ;
        RECT -16.220 1476.990 -15.040 1478.170 ;
        RECT -14.620 1476.990 -13.440 1478.170 ;
        RECT -16.220 1298.590 -15.040 1299.770 ;
        RECT -14.620 1298.590 -13.440 1299.770 ;
        RECT -16.220 1296.990 -15.040 1298.170 ;
        RECT -14.620 1296.990 -13.440 1298.170 ;
        RECT -16.220 1118.590 -15.040 1119.770 ;
        RECT -14.620 1118.590 -13.440 1119.770 ;
        RECT -16.220 1116.990 -15.040 1118.170 ;
        RECT -14.620 1116.990 -13.440 1118.170 ;
        RECT -16.220 938.590 -15.040 939.770 ;
        RECT -14.620 938.590 -13.440 939.770 ;
        RECT -16.220 936.990 -15.040 938.170 ;
        RECT -14.620 936.990 -13.440 938.170 ;
        RECT -16.220 758.590 -15.040 759.770 ;
        RECT -14.620 758.590 -13.440 759.770 ;
        RECT -16.220 756.990 -15.040 758.170 ;
        RECT -14.620 756.990 -13.440 758.170 ;
        RECT -16.220 578.590 -15.040 579.770 ;
        RECT -14.620 578.590 -13.440 579.770 ;
        RECT -16.220 576.990 -15.040 578.170 ;
        RECT -14.620 576.990 -13.440 578.170 ;
        RECT -16.220 398.590 -15.040 399.770 ;
        RECT -14.620 398.590 -13.440 399.770 ;
        RECT -16.220 396.990 -15.040 398.170 ;
        RECT -14.620 396.990 -13.440 398.170 ;
        RECT -16.220 218.590 -15.040 219.770 ;
        RECT -14.620 218.590 -13.440 219.770 ;
        RECT -16.220 216.990 -15.040 218.170 ;
        RECT -14.620 216.990 -13.440 218.170 ;
        RECT -16.220 38.590 -15.040 39.770 ;
        RECT -14.620 38.590 -13.440 39.770 ;
        RECT -16.220 36.990 -15.040 38.170 ;
        RECT -14.620 36.990 -13.440 38.170 ;
        RECT -16.220 -9.260 -15.040 -8.080 ;
        RECT -14.620 -9.260 -13.440 -8.080 ;
        RECT -16.220 -10.860 -15.040 -9.680 ;
        RECT -14.620 -10.860 -13.440 -9.680 ;
        RECT 31.630 3529.360 32.810 3530.540 ;
        RECT 33.230 3529.360 34.410 3530.540 ;
        RECT 31.630 3527.760 32.810 3528.940 ;
        RECT 33.230 3527.760 34.410 3528.940 ;
        RECT 31.630 3458.590 32.810 3459.770 ;
        RECT 33.230 3458.590 34.410 3459.770 ;
        RECT 31.630 3456.990 32.810 3458.170 ;
        RECT 33.230 3456.990 34.410 3458.170 ;
        RECT 31.630 3278.590 32.810 3279.770 ;
        RECT 33.230 3278.590 34.410 3279.770 ;
        RECT 31.630 3276.990 32.810 3278.170 ;
        RECT 33.230 3276.990 34.410 3278.170 ;
        RECT 31.630 3098.590 32.810 3099.770 ;
        RECT 33.230 3098.590 34.410 3099.770 ;
        RECT 31.630 3096.990 32.810 3098.170 ;
        RECT 33.230 3096.990 34.410 3098.170 ;
        RECT 31.630 2918.590 32.810 2919.770 ;
        RECT 33.230 2918.590 34.410 2919.770 ;
        RECT 31.630 2916.990 32.810 2918.170 ;
        RECT 33.230 2916.990 34.410 2918.170 ;
        RECT 31.630 2738.590 32.810 2739.770 ;
        RECT 33.230 2738.590 34.410 2739.770 ;
        RECT 31.630 2736.990 32.810 2738.170 ;
        RECT 33.230 2736.990 34.410 2738.170 ;
        RECT 31.630 2558.590 32.810 2559.770 ;
        RECT 33.230 2558.590 34.410 2559.770 ;
        RECT 31.630 2556.990 32.810 2558.170 ;
        RECT 33.230 2556.990 34.410 2558.170 ;
        RECT 31.630 2378.590 32.810 2379.770 ;
        RECT 33.230 2378.590 34.410 2379.770 ;
        RECT 31.630 2376.990 32.810 2378.170 ;
        RECT 33.230 2376.990 34.410 2378.170 ;
        RECT 31.630 2198.590 32.810 2199.770 ;
        RECT 33.230 2198.590 34.410 2199.770 ;
        RECT 31.630 2196.990 32.810 2198.170 ;
        RECT 33.230 2196.990 34.410 2198.170 ;
        RECT 31.630 2018.590 32.810 2019.770 ;
        RECT 33.230 2018.590 34.410 2019.770 ;
        RECT 31.630 2016.990 32.810 2018.170 ;
        RECT 33.230 2016.990 34.410 2018.170 ;
        RECT 31.630 1838.590 32.810 1839.770 ;
        RECT 33.230 1838.590 34.410 1839.770 ;
        RECT 31.630 1836.990 32.810 1838.170 ;
        RECT 33.230 1836.990 34.410 1838.170 ;
        RECT 31.630 1658.590 32.810 1659.770 ;
        RECT 33.230 1658.590 34.410 1659.770 ;
        RECT 31.630 1656.990 32.810 1658.170 ;
        RECT 33.230 1656.990 34.410 1658.170 ;
        RECT 31.630 1478.590 32.810 1479.770 ;
        RECT 33.230 1478.590 34.410 1479.770 ;
        RECT 31.630 1476.990 32.810 1478.170 ;
        RECT 33.230 1476.990 34.410 1478.170 ;
        RECT 31.630 1298.590 32.810 1299.770 ;
        RECT 33.230 1298.590 34.410 1299.770 ;
        RECT 31.630 1296.990 32.810 1298.170 ;
        RECT 33.230 1296.990 34.410 1298.170 ;
        RECT 31.630 1118.590 32.810 1119.770 ;
        RECT 33.230 1118.590 34.410 1119.770 ;
        RECT 31.630 1116.990 32.810 1118.170 ;
        RECT 33.230 1116.990 34.410 1118.170 ;
        RECT 31.630 938.590 32.810 939.770 ;
        RECT 33.230 938.590 34.410 939.770 ;
        RECT 31.630 936.990 32.810 938.170 ;
        RECT 33.230 936.990 34.410 938.170 ;
        RECT 31.630 758.590 32.810 759.770 ;
        RECT 33.230 758.590 34.410 759.770 ;
        RECT 31.630 756.990 32.810 758.170 ;
        RECT 33.230 756.990 34.410 758.170 ;
        RECT 31.630 578.590 32.810 579.770 ;
        RECT 33.230 578.590 34.410 579.770 ;
        RECT 31.630 576.990 32.810 578.170 ;
        RECT 33.230 576.990 34.410 578.170 ;
        RECT 31.630 398.590 32.810 399.770 ;
        RECT 33.230 398.590 34.410 399.770 ;
        RECT 31.630 396.990 32.810 398.170 ;
        RECT 33.230 396.990 34.410 398.170 ;
        RECT 31.630 218.590 32.810 219.770 ;
        RECT 33.230 218.590 34.410 219.770 ;
        RECT 31.630 216.990 32.810 218.170 ;
        RECT 33.230 216.990 34.410 218.170 ;
        RECT 31.630 38.590 32.810 39.770 ;
        RECT 33.230 38.590 34.410 39.770 ;
        RECT 31.630 36.990 32.810 38.170 ;
        RECT 33.230 36.990 34.410 38.170 ;
        RECT 31.630 -9.260 32.810 -8.080 ;
        RECT 33.230 -9.260 34.410 -8.080 ;
        RECT 31.630 -10.860 32.810 -9.680 ;
        RECT 33.230 -10.860 34.410 -9.680 ;
        RECT 211.630 3529.360 212.810 3530.540 ;
        RECT 213.230 3529.360 214.410 3530.540 ;
        RECT 211.630 3527.760 212.810 3528.940 ;
        RECT 213.230 3527.760 214.410 3528.940 ;
        RECT 211.630 3458.590 212.810 3459.770 ;
        RECT 213.230 3458.590 214.410 3459.770 ;
        RECT 211.630 3456.990 212.810 3458.170 ;
        RECT 213.230 3456.990 214.410 3458.170 ;
        RECT 211.630 3278.590 212.810 3279.770 ;
        RECT 213.230 3278.590 214.410 3279.770 ;
        RECT 211.630 3276.990 212.810 3278.170 ;
        RECT 213.230 3276.990 214.410 3278.170 ;
        RECT 211.630 3098.590 212.810 3099.770 ;
        RECT 213.230 3098.590 214.410 3099.770 ;
        RECT 211.630 3096.990 212.810 3098.170 ;
        RECT 213.230 3096.990 214.410 3098.170 ;
        RECT 211.630 2918.590 212.810 2919.770 ;
        RECT 213.230 2918.590 214.410 2919.770 ;
        RECT 211.630 2916.990 212.810 2918.170 ;
        RECT 213.230 2916.990 214.410 2918.170 ;
        RECT 211.630 2738.590 212.810 2739.770 ;
        RECT 213.230 2738.590 214.410 2739.770 ;
        RECT 211.630 2736.990 212.810 2738.170 ;
        RECT 213.230 2736.990 214.410 2738.170 ;
        RECT 211.630 2558.590 212.810 2559.770 ;
        RECT 213.230 2558.590 214.410 2559.770 ;
        RECT 211.630 2556.990 212.810 2558.170 ;
        RECT 213.230 2556.990 214.410 2558.170 ;
        RECT 211.630 2378.590 212.810 2379.770 ;
        RECT 213.230 2378.590 214.410 2379.770 ;
        RECT 211.630 2376.990 212.810 2378.170 ;
        RECT 213.230 2376.990 214.410 2378.170 ;
        RECT 211.630 2198.590 212.810 2199.770 ;
        RECT 213.230 2198.590 214.410 2199.770 ;
        RECT 211.630 2196.990 212.810 2198.170 ;
        RECT 213.230 2196.990 214.410 2198.170 ;
        RECT 211.630 2018.590 212.810 2019.770 ;
        RECT 213.230 2018.590 214.410 2019.770 ;
        RECT 211.630 2016.990 212.810 2018.170 ;
        RECT 213.230 2016.990 214.410 2018.170 ;
        RECT 211.630 1838.590 212.810 1839.770 ;
        RECT 213.230 1838.590 214.410 1839.770 ;
        RECT 211.630 1836.990 212.810 1838.170 ;
        RECT 213.230 1836.990 214.410 1838.170 ;
        RECT 211.630 1658.590 212.810 1659.770 ;
        RECT 213.230 1658.590 214.410 1659.770 ;
        RECT 211.630 1656.990 212.810 1658.170 ;
        RECT 213.230 1656.990 214.410 1658.170 ;
        RECT 211.630 1478.590 212.810 1479.770 ;
        RECT 213.230 1478.590 214.410 1479.770 ;
        RECT 211.630 1476.990 212.810 1478.170 ;
        RECT 213.230 1476.990 214.410 1478.170 ;
        RECT 211.630 1298.590 212.810 1299.770 ;
        RECT 213.230 1298.590 214.410 1299.770 ;
        RECT 211.630 1296.990 212.810 1298.170 ;
        RECT 213.230 1296.990 214.410 1298.170 ;
        RECT 211.630 1118.590 212.810 1119.770 ;
        RECT 213.230 1118.590 214.410 1119.770 ;
        RECT 211.630 1116.990 212.810 1118.170 ;
        RECT 213.230 1116.990 214.410 1118.170 ;
        RECT 211.630 938.590 212.810 939.770 ;
        RECT 213.230 938.590 214.410 939.770 ;
        RECT 211.630 936.990 212.810 938.170 ;
        RECT 213.230 936.990 214.410 938.170 ;
        RECT 391.630 3529.360 392.810 3530.540 ;
        RECT 393.230 3529.360 394.410 3530.540 ;
        RECT 391.630 3527.760 392.810 3528.940 ;
        RECT 393.230 3527.760 394.410 3528.940 ;
        RECT 391.630 3458.590 392.810 3459.770 ;
        RECT 393.230 3458.590 394.410 3459.770 ;
        RECT 391.630 3456.990 392.810 3458.170 ;
        RECT 393.230 3456.990 394.410 3458.170 ;
        RECT 391.630 3278.590 392.810 3279.770 ;
        RECT 393.230 3278.590 394.410 3279.770 ;
        RECT 391.630 3276.990 392.810 3278.170 ;
        RECT 393.230 3276.990 394.410 3278.170 ;
        RECT 391.630 3098.590 392.810 3099.770 ;
        RECT 393.230 3098.590 394.410 3099.770 ;
        RECT 391.630 3096.990 392.810 3098.170 ;
        RECT 393.230 3096.990 394.410 3098.170 ;
        RECT 391.630 2918.590 392.810 2919.770 ;
        RECT 393.230 2918.590 394.410 2919.770 ;
        RECT 391.630 2916.990 392.810 2918.170 ;
        RECT 393.230 2916.990 394.410 2918.170 ;
        RECT 391.630 2738.590 392.810 2739.770 ;
        RECT 393.230 2738.590 394.410 2739.770 ;
        RECT 391.630 2736.990 392.810 2738.170 ;
        RECT 393.230 2736.990 394.410 2738.170 ;
        RECT 391.630 2558.590 392.810 2559.770 ;
        RECT 393.230 2558.590 394.410 2559.770 ;
        RECT 391.630 2556.990 392.810 2558.170 ;
        RECT 393.230 2556.990 394.410 2558.170 ;
        RECT 391.630 2378.590 392.810 2379.770 ;
        RECT 393.230 2378.590 394.410 2379.770 ;
        RECT 391.630 2376.990 392.810 2378.170 ;
        RECT 393.230 2376.990 394.410 2378.170 ;
        RECT 391.630 2198.590 392.810 2199.770 ;
        RECT 393.230 2198.590 394.410 2199.770 ;
        RECT 391.630 2196.990 392.810 2198.170 ;
        RECT 393.230 2196.990 394.410 2198.170 ;
        RECT 391.630 2018.590 392.810 2019.770 ;
        RECT 393.230 2018.590 394.410 2019.770 ;
        RECT 391.630 2016.990 392.810 2018.170 ;
        RECT 393.230 2016.990 394.410 2018.170 ;
        RECT 391.630 1838.590 392.810 1839.770 ;
        RECT 393.230 1838.590 394.410 1839.770 ;
        RECT 391.630 1836.990 392.810 1838.170 ;
        RECT 393.230 1836.990 394.410 1838.170 ;
        RECT 391.630 1658.590 392.810 1659.770 ;
        RECT 393.230 1658.590 394.410 1659.770 ;
        RECT 391.630 1656.990 392.810 1658.170 ;
        RECT 393.230 1656.990 394.410 1658.170 ;
        RECT 391.630 1478.590 392.810 1479.770 ;
        RECT 393.230 1478.590 394.410 1479.770 ;
        RECT 391.630 1476.990 392.810 1478.170 ;
        RECT 393.230 1476.990 394.410 1478.170 ;
        RECT 391.630 1298.590 392.810 1299.770 ;
        RECT 393.230 1298.590 394.410 1299.770 ;
        RECT 391.630 1296.990 392.810 1298.170 ;
        RECT 393.230 1296.990 394.410 1298.170 ;
        RECT 391.630 1118.590 392.810 1119.770 ;
        RECT 393.230 1118.590 394.410 1119.770 ;
        RECT 391.630 1116.990 392.810 1118.170 ;
        RECT 393.230 1116.990 394.410 1118.170 ;
        RECT 391.630 938.590 392.810 939.770 ;
        RECT 393.230 938.590 394.410 939.770 ;
        RECT 391.630 936.990 392.810 938.170 ;
        RECT 393.230 936.990 394.410 938.170 ;
        RECT 571.630 3529.360 572.810 3530.540 ;
        RECT 573.230 3529.360 574.410 3530.540 ;
        RECT 571.630 3527.760 572.810 3528.940 ;
        RECT 573.230 3527.760 574.410 3528.940 ;
        RECT 571.630 3458.590 572.810 3459.770 ;
        RECT 573.230 3458.590 574.410 3459.770 ;
        RECT 571.630 3456.990 572.810 3458.170 ;
        RECT 573.230 3456.990 574.410 3458.170 ;
        RECT 571.630 3278.590 572.810 3279.770 ;
        RECT 573.230 3278.590 574.410 3279.770 ;
        RECT 571.630 3276.990 572.810 3278.170 ;
        RECT 573.230 3276.990 574.410 3278.170 ;
        RECT 571.630 3098.590 572.810 3099.770 ;
        RECT 573.230 3098.590 574.410 3099.770 ;
        RECT 571.630 3096.990 572.810 3098.170 ;
        RECT 573.230 3096.990 574.410 3098.170 ;
        RECT 571.630 2918.590 572.810 2919.770 ;
        RECT 573.230 2918.590 574.410 2919.770 ;
        RECT 571.630 2916.990 572.810 2918.170 ;
        RECT 573.230 2916.990 574.410 2918.170 ;
        RECT 571.630 2738.590 572.810 2739.770 ;
        RECT 573.230 2738.590 574.410 2739.770 ;
        RECT 571.630 2736.990 572.810 2738.170 ;
        RECT 573.230 2736.990 574.410 2738.170 ;
        RECT 571.630 2558.590 572.810 2559.770 ;
        RECT 573.230 2558.590 574.410 2559.770 ;
        RECT 571.630 2556.990 572.810 2558.170 ;
        RECT 573.230 2556.990 574.410 2558.170 ;
        RECT 571.630 2378.590 572.810 2379.770 ;
        RECT 573.230 2378.590 574.410 2379.770 ;
        RECT 571.630 2376.990 572.810 2378.170 ;
        RECT 573.230 2376.990 574.410 2378.170 ;
        RECT 571.630 2198.590 572.810 2199.770 ;
        RECT 573.230 2198.590 574.410 2199.770 ;
        RECT 571.630 2196.990 572.810 2198.170 ;
        RECT 573.230 2196.990 574.410 2198.170 ;
        RECT 571.630 2018.590 572.810 2019.770 ;
        RECT 573.230 2018.590 574.410 2019.770 ;
        RECT 571.630 2016.990 572.810 2018.170 ;
        RECT 573.230 2016.990 574.410 2018.170 ;
        RECT 571.630 1838.590 572.810 1839.770 ;
        RECT 573.230 1838.590 574.410 1839.770 ;
        RECT 571.630 1836.990 572.810 1838.170 ;
        RECT 573.230 1836.990 574.410 1838.170 ;
        RECT 571.630 1658.590 572.810 1659.770 ;
        RECT 573.230 1658.590 574.410 1659.770 ;
        RECT 571.630 1656.990 572.810 1658.170 ;
        RECT 573.230 1656.990 574.410 1658.170 ;
        RECT 571.630 1478.590 572.810 1479.770 ;
        RECT 573.230 1478.590 574.410 1479.770 ;
        RECT 571.630 1476.990 572.810 1478.170 ;
        RECT 573.230 1476.990 574.410 1478.170 ;
        RECT 571.630 1298.590 572.810 1299.770 ;
        RECT 573.230 1298.590 574.410 1299.770 ;
        RECT 571.630 1296.990 572.810 1298.170 ;
        RECT 573.230 1296.990 574.410 1298.170 ;
        RECT 571.630 1118.590 572.810 1119.770 ;
        RECT 573.230 1118.590 574.410 1119.770 ;
        RECT 571.630 1116.990 572.810 1118.170 ;
        RECT 573.230 1116.990 574.410 1118.170 ;
        RECT 571.630 938.590 572.810 939.770 ;
        RECT 573.230 938.590 574.410 939.770 ;
        RECT 571.630 936.990 572.810 938.170 ;
        RECT 573.230 936.990 574.410 938.170 ;
        RECT 751.630 3529.360 752.810 3530.540 ;
        RECT 753.230 3529.360 754.410 3530.540 ;
        RECT 751.630 3527.760 752.810 3528.940 ;
        RECT 753.230 3527.760 754.410 3528.940 ;
        RECT 751.630 3458.590 752.810 3459.770 ;
        RECT 753.230 3458.590 754.410 3459.770 ;
        RECT 751.630 3456.990 752.810 3458.170 ;
        RECT 753.230 3456.990 754.410 3458.170 ;
        RECT 751.630 3278.590 752.810 3279.770 ;
        RECT 753.230 3278.590 754.410 3279.770 ;
        RECT 751.630 3276.990 752.810 3278.170 ;
        RECT 753.230 3276.990 754.410 3278.170 ;
        RECT 751.630 3098.590 752.810 3099.770 ;
        RECT 753.230 3098.590 754.410 3099.770 ;
        RECT 751.630 3096.990 752.810 3098.170 ;
        RECT 753.230 3096.990 754.410 3098.170 ;
        RECT 751.630 2918.590 752.810 2919.770 ;
        RECT 753.230 2918.590 754.410 2919.770 ;
        RECT 751.630 2916.990 752.810 2918.170 ;
        RECT 753.230 2916.990 754.410 2918.170 ;
        RECT 751.630 2738.590 752.810 2739.770 ;
        RECT 753.230 2738.590 754.410 2739.770 ;
        RECT 751.630 2736.990 752.810 2738.170 ;
        RECT 753.230 2736.990 754.410 2738.170 ;
        RECT 751.630 2558.590 752.810 2559.770 ;
        RECT 753.230 2558.590 754.410 2559.770 ;
        RECT 751.630 2556.990 752.810 2558.170 ;
        RECT 753.230 2556.990 754.410 2558.170 ;
        RECT 751.630 2378.590 752.810 2379.770 ;
        RECT 753.230 2378.590 754.410 2379.770 ;
        RECT 751.630 2376.990 752.810 2378.170 ;
        RECT 753.230 2376.990 754.410 2378.170 ;
        RECT 751.630 2198.590 752.810 2199.770 ;
        RECT 753.230 2198.590 754.410 2199.770 ;
        RECT 751.630 2196.990 752.810 2198.170 ;
        RECT 753.230 2196.990 754.410 2198.170 ;
        RECT 751.630 2018.590 752.810 2019.770 ;
        RECT 753.230 2018.590 754.410 2019.770 ;
        RECT 751.630 2016.990 752.810 2018.170 ;
        RECT 753.230 2016.990 754.410 2018.170 ;
        RECT 751.630 1838.590 752.810 1839.770 ;
        RECT 753.230 1838.590 754.410 1839.770 ;
        RECT 751.630 1836.990 752.810 1838.170 ;
        RECT 753.230 1836.990 754.410 1838.170 ;
        RECT 751.630 1658.590 752.810 1659.770 ;
        RECT 753.230 1658.590 754.410 1659.770 ;
        RECT 751.630 1656.990 752.810 1658.170 ;
        RECT 753.230 1656.990 754.410 1658.170 ;
        RECT 751.630 1478.590 752.810 1479.770 ;
        RECT 753.230 1478.590 754.410 1479.770 ;
        RECT 751.630 1476.990 752.810 1478.170 ;
        RECT 753.230 1476.990 754.410 1478.170 ;
        RECT 751.630 1298.590 752.810 1299.770 ;
        RECT 753.230 1298.590 754.410 1299.770 ;
        RECT 751.630 1296.990 752.810 1298.170 ;
        RECT 753.230 1296.990 754.410 1298.170 ;
        RECT 751.630 1118.590 752.810 1119.770 ;
        RECT 753.230 1118.590 754.410 1119.770 ;
        RECT 751.630 1116.990 752.810 1118.170 ;
        RECT 753.230 1116.990 754.410 1118.170 ;
        RECT 751.630 938.590 752.810 939.770 ;
        RECT 753.230 938.590 754.410 939.770 ;
        RECT 751.630 936.990 752.810 938.170 ;
        RECT 753.230 936.990 754.410 938.170 ;
        RECT 211.630 758.590 212.810 759.770 ;
        RECT 213.230 758.590 214.410 759.770 ;
        RECT 211.630 756.990 212.810 758.170 ;
        RECT 213.230 756.990 214.410 758.170 ;
        RECT 751.630 758.590 752.810 759.770 ;
        RECT 753.230 758.590 754.410 759.770 ;
        RECT 751.630 756.990 752.810 758.170 ;
        RECT 753.230 756.990 754.410 758.170 ;
        RECT 211.630 578.590 212.810 579.770 ;
        RECT 213.230 578.590 214.410 579.770 ;
        RECT 211.630 576.990 212.810 578.170 ;
        RECT 213.230 576.990 214.410 578.170 ;
        RECT 498.050 578.590 499.230 579.770 ;
        RECT 498.050 576.990 499.230 578.170 ;
        RECT 751.630 578.590 752.810 579.770 ;
        RECT 753.230 578.590 754.410 579.770 ;
        RECT 751.630 576.990 752.810 578.170 ;
        RECT 753.230 576.990 754.410 578.170 ;
        RECT 211.630 398.590 212.810 399.770 ;
        RECT 213.230 398.590 214.410 399.770 ;
        RECT 211.630 396.990 212.810 398.170 ;
        RECT 213.230 396.990 214.410 398.170 ;
        RECT 211.630 218.590 212.810 219.770 ;
        RECT 213.230 218.590 214.410 219.770 ;
        RECT 211.630 216.990 212.810 218.170 ;
        RECT 213.230 216.990 214.410 218.170 ;
        RECT 211.630 38.590 212.810 39.770 ;
        RECT 213.230 38.590 214.410 39.770 ;
        RECT 211.630 36.990 212.810 38.170 ;
        RECT 213.230 36.990 214.410 38.170 ;
        RECT 211.630 -9.260 212.810 -8.080 ;
        RECT 213.230 -9.260 214.410 -8.080 ;
        RECT 211.630 -10.860 212.810 -9.680 ;
        RECT 213.230 -10.860 214.410 -9.680 ;
        RECT 391.630 398.590 392.810 399.770 ;
        RECT 393.230 398.590 394.410 399.770 ;
        RECT 391.630 396.990 392.810 398.170 ;
        RECT 393.230 396.990 394.410 398.170 ;
        RECT 391.630 218.590 392.810 219.770 ;
        RECT 393.230 218.590 394.410 219.770 ;
        RECT 391.630 216.990 392.810 218.170 ;
        RECT 393.230 216.990 394.410 218.170 ;
        RECT 391.630 38.590 392.810 39.770 ;
        RECT 393.230 38.590 394.410 39.770 ;
        RECT 391.630 36.990 392.810 38.170 ;
        RECT 393.230 36.990 394.410 38.170 ;
        RECT 391.630 -9.260 392.810 -8.080 ;
        RECT 393.230 -9.260 394.410 -8.080 ;
        RECT 391.630 -10.860 392.810 -9.680 ;
        RECT 393.230 -10.860 394.410 -9.680 ;
        RECT 571.630 398.590 572.810 399.770 ;
        RECT 573.230 398.590 574.410 399.770 ;
        RECT 571.630 396.990 572.810 398.170 ;
        RECT 573.230 396.990 574.410 398.170 ;
        RECT 571.630 218.590 572.810 219.770 ;
        RECT 573.230 218.590 574.410 219.770 ;
        RECT 571.630 216.990 572.810 218.170 ;
        RECT 573.230 216.990 574.410 218.170 ;
        RECT 571.630 38.590 572.810 39.770 ;
        RECT 573.230 38.590 574.410 39.770 ;
        RECT 571.630 36.990 572.810 38.170 ;
        RECT 573.230 36.990 574.410 38.170 ;
        RECT 571.630 -9.260 572.810 -8.080 ;
        RECT 573.230 -9.260 574.410 -8.080 ;
        RECT 571.630 -10.860 572.810 -9.680 ;
        RECT 573.230 -10.860 574.410 -9.680 ;
        RECT 751.630 398.590 752.810 399.770 ;
        RECT 753.230 398.590 754.410 399.770 ;
        RECT 751.630 396.990 752.810 398.170 ;
        RECT 753.230 396.990 754.410 398.170 ;
        RECT 751.630 218.590 752.810 219.770 ;
        RECT 753.230 218.590 754.410 219.770 ;
        RECT 751.630 216.990 752.810 218.170 ;
        RECT 753.230 216.990 754.410 218.170 ;
        RECT 751.630 38.590 752.810 39.770 ;
        RECT 753.230 38.590 754.410 39.770 ;
        RECT 751.630 36.990 752.810 38.170 ;
        RECT 753.230 36.990 754.410 38.170 ;
        RECT 751.630 -9.260 752.810 -8.080 ;
        RECT 753.230 -9.260 754.410 -8.080 ;
        RECT 751.630 -10.860 752.810 -9.680 ;
        RECT 753.230 -10.860 754.410 -9.680 ;
        RECT 931.630 3529.360 932.810 3530.540 ;
        RECT 933.230 3529.360 934.410 3530.540 ;
        RECT 931.630 3527.760 932.810 3528.940 ;
        RECT 933.230 3527.760 934.410 3528.940 ;
        RECT 931.630 3458.590 932.810 3459.770 ;
        RECT 933.230 3458.590 934.410 3459.770 ;
        RECT 931.630 3456.990 932.810 3458.170 ;
        RECT 933.230 3456.990 934.410 3458.170 ;
        RECT 931.630 3278.590 932.810 3279.770 ;
        RECT 933.230 3278.590 934.410 3279.770 ;
        RECT 931.630 3276.990 932.810 3278.170 ;
        RECT 933.230 3276.990 934.410 3278.170 ;
        RECT 931.630 3098.590 932.810 3099.770 ;
        RECT 933.230 3098.590 934.410 3099.770 ;
        RECT 931.630 3096.990 932.810 3098.170 ;
        RECT 933.230 3096.990 934.410 3098.170 ;
        RECT 931.630 2918.590 932.810 2919.770 ;
        RECT 933.230 2918.590 934.410 2919.770 ;
        RECT 931.630 2916.990 932.810 2918.170 ;
        RECT 933.230 2916.990 934.410 2918.170 ;
        RECT 931.630 2738.590 932.810 2739.770 ;
        RECT 933.230 2738.590 934.410 2739.770 ;
        RECT 931.630 2736.990 932.810 2738.170 ;
        RECT 933.230 2736.990 934.410 2738.170 ;
        RECT 931.630 2558.590 932.810 2559.770 ;
        RECT 933.230 2558.590 934.410 2559.770 ;
        RECT 931.630 2556.990 932.810 2558.170 ;
        RECT 933.230 2556.990 934.410 2558.170 ;
        RECT 931.630 2378.590 932.810 2379.770 ;
        RECT 933.230 2378.590 934.410 2379.770 ;
        RECT 931.630 2376.990 932.810 2378.170 ;
        RECT 933.230 2376.990 934.410 2378.170 ;
        RECT 931.630 2198.590 932.810 2199.770 ;
        RECT 933.230 2198.590 934.410 2199.770 ;
        RECT 931.630 2196.990 932.810 2198.170 ;
        RECT 933.230 2196.990 934.410 2198.170 ;
        RECT 931.630 2018.590 932.810 2019.770 ;
        RECT 933.230 2018.590 934.410 2019.770 ;
        RECT 931.630 2016.990 932.810 2018.170 ;
        RECT 933.230 2016.990 934.410 2018.170 ;
        RECT 931.630 1838.590 932.810 1839.770 ;
        RECT 933.230 1838.590 934.410 1839.770 ;
        RECT 931.630 1836.990 932.810 1838.170 ;
        RECT 933.230 1836.990 934.410 1838.170 ;
        RECT 931.630 1658.590 932.810 1659.770 ;
        RECT 933.230 1658.590 934.410 1659.770 ;
        RECT 931.630 1656.990 932.810 1658.170 ;
        RECT 933.230 1656.990 934.410 1658.170 ;
        RECT 931.630 1478.590 932.810 1479.770 ;
        RECT 933.230 1478.590 934.410 1479.770 ;
        RECT 931.630 1476.990 932.810 1478.170 ;
        RECT 933.230 1476.990 934.410 1478.170 ;
        RECT 931.630 1298.590 932.810 1299.770 ;
        RECT 933.230 1298.590 934.410 1299.770 ;
        RECT 931.630 1296.990 932.810 1298.170 ;
        RECT 933.230 1296.990 934.410 1298.170 ;
        RECT 931.630 1118.590 932.810 1119.770 ;
        RECT 933.230 1118.590 934.410 1119.770 ;
        RECT 931.630 1116.990 932.810 1118.170 ;
        RECT 933.230 1116.990 934.410 1118.170 ;
        RECT 931.630 938.590 932.810 939.770 ;
        RECT 933.230 938.590 934.410 939.770 ;
        RECT 931.630 936.990 932.810 938.170 ;
        RECT 933.230 936.990 934.410 938.170 ;
        RECT 931.630 758.590 932.810 759.770 ;
        RECT 933.230 758.590 934.410 759.770 ;
        RECT 931.630 756.990 932.810 758.170 ;
        RECT 933.230 756.990 934.410 758.170 ;
        RECT 931.630 578.590 932.810 579.770 ;
        RECT 933.230 578.590 934.410 579.770 ;
        RECT 931.630 576.990 932.810 578.170 ;
        RECT 933.230 576.990 934.410 578.170 ;
        RECT 931.630 398.590 932.810 399.770 ;
        RECT 933.230 398.590 934.410 399.770 ;
        RECT 931.630 396.990 932.810 398.170 ;
        RECT 933.230 396.990 934.410 398.170 ;
        RECT 931.630 218.590 932.810 219.770 ;
        RECT 933.230 218.590 934.410 219.770 ;
        RECT 931.630 216.990 932.810 218.170 ;
        RECT 933.230 216.990 934.410 218.170 ;
        RECT 931.630 38.590 932.810 39.770 ;
        RECT 933.230 38.590 934.410 39.770 ;
        RECT 931.630 36.990 932.810 38.170 ;
        RECT 933.230 36.990 934.410 38.170 ;
        RECT 931.630 -9.260 932.810 -8.080 ;
        RECT 933.230 -9.260 934.410 -8.080 ;
        RECT 931.630 -10.860 932.810 -9.680 ;
        RECT 933.230 -10.860 934.410 -9.680 ;
        RECT 1111.630 3529.360 1112.810 3530.540 ;
        RECT 1113.230 3529.360 1114.410 3530.540 ;
        RECT 1111.630 3527.760 1112.810 3528.940 ;
        RECT 1113.230 3527.760 1114.410 3528.940 ;
        RECT 1111.630 3458.590 1112.810 3459.770 ;
        RECT 1113.230 3458.590 1114.410 3459.770 ;
        RECT 1111.630 3456.990 1112.810 3458.170 ;
        RECT 1113.230 3456.990 1114.410 3458.170 ;
        RECT 1111.630 3278.590 1112.810 3279.770 ;
        RECT 1113.230 3278.590 1114.410 3279.770 ;
        RECT 1111.630 3276.990 1112.810 3278.170 ;
        RECT 1113.230 3276.990 1114.410 3278.170 ;
        RECT 1111.630 3098.590 1112.810 3099.770 ;
        RECT 1113.230 3098.590 1114.410 3099.770 ;
        RECT 1111.630 3096.990 1112.810 3098.170 ;
        RECT 1113.230 3096.990 1114.410 3098.170 ;
        RECT 1111.630 2918.590 1112.810 2919.770 ;
        RECT 1113.230 2918.590 1114.410 2919.770 ;
        RECT 1111.630 2916.990 1112.810 2918.170 ;
        RECT 1113.230 2916.990 1114.410 2918.170 ;
        RECT 1111.630 2738.590 1112.810 2739.770 ;
        RECT 1113.230 2738.590 1114.410 2739.770 ;
        RECT 1111.630 2736.990 1112.810 2738.170 ;
        RECT 1113.230 2736.990 1114.410 2738.170 ;
        RECT 1111.630 2558.590 1112.810 2559.770 ;
        RECT 1113.230 2558.590 1114.410 2559.770 ;
        RECT 1111.630 2556.990 1112.810 2558.170 ;
        RECT 1113.230 2556.990 1114.410 2558.170 ;
        RECT 1111.630 2378.590 1112.810 2379.770 ;
        RECT 1113.230 2378.590 1114.410 2379.770 ;
        RECT 1111.630 2376.990 1112.810 2378.170 ;
        RECT 1113.230 2376.990 1114.410 2378.170 ;
        RECT 1111.630 2198.590 1112.810 2199.770 ;
        RECT 1113.230 2198.590 1114.410 2199.770 ;
        RECT 1111.630 2196.990 1112.810 2198.170 ;
        RECT 1113.230 2196.990 1114.410 2198.170 ;
        RECT 1111.630 2018.590 1112.810 2019.770 ;
        RECT 1113.230 2018.590 1114.410 2019.770 ;
        RECT 1111.630 2016.990 1112.810 2018.170 ;
        RECT 1113.230 2016.990 1114.410 2018.170 ;
        RECT 1111.630 1838.590 1112.810 1839.770 ;
        RECT 1113.230 1838.590 1114.410 1839.770 ;
        RECT 1111.630 1836.990 1112.810 1838.170 ;
        RECT 1113.230 1836.990 1114.410 1838.170 ;
        RECT 1111.630 1658.590 1112.810 1659.770 ;
        RECT 1113.230 1658.590 1114.410 1659.770 ;
        RECT 1111.630 1656.990 1112.810 1658.170 ;
        RECT 1113.230 1656.990 1114.410 1658.170 ;
        RECT 1111.630 1478.590 1112.810 1479.770 ;
        RECT 1113.230 1478.590 1114.410 1479.770 ;
        RECT 1111.630 1476.990 1112.810 1478.170 ;
        RECT 1113.230 1476.990 1114.410 1478.170 ;
        RECT 1111.630 1298.590 1112.810 1299.770 ;
        RECT 1113.230 1298.590 1114.410 1299.770 ;
        RECT 1111.630 1296.990 1112.810 1298.170 ;
        RECT 1113.230 1296.990 1114.410 1298.170 ;
        RECT 1111.630 1118.590 1112.810 1119.770 ;
        RECT 1113.230 1118.590 1114.410 1119.770 ;
        RECT 1111.630 1116.990 1112.810 1118.170 ;
        RECT 1113.230 1116.990 1114.410 1118.170 ;
        RECT 1111.630 938.590 1112.810 939.770 ;
        RECT 1113.230 938.590 1114.410 939.770 ;
        RECT 1111.630 936.990 1112.810 938.170 ;
        RECT 1113.230 936.990 1114.410 938.170 ;
        RECT 1111.630 758.590 1112.810 759.770 ;
        RECT 1113.230 758.590 1114.410 759.770 ;
        RECT 1111.630 756.990 1112.810 758.170 ;
        RECT 1113.230 756.990 1114.410 758.170 ;
        RECT 1111.630 578.590 1112.810 579.770 ;
        RECT 1113.230 578.590 1114.410 579.770 ;
        RECT 1111.630 576.990 1112.810 578.170 ;
        RECT 1113.230 576.990 1114.410 578.170 ;
        RECT 1111.630 398.590 1112.810 399.770 ;
        RECT 1113.230 398.590 1114.410 399.770 ;
        RECT 1111.630 396.990 1112.810 398.170 ;
        RECT 1113.230 396.990 1114.410 398.170 ;
        RECT 1111.630 218.590 1112.810 219.770 ;
        RECT 1113.230 218.590 1114.410 219.770 ;
        RECT 1111.630 216.990 1112.810 218.170 ;
        RECT 1113.230 216.990 1114.410 218.170 ;
        RECT 1111.630 38.590 1112.810 39.770 ;
        RECT 1113.230 38.590 1114.410 39.770 ;
        RECT 1111.630 36.990 1112.810 38.170 ;
        RECT 1113.230 36.990 1114.410 38.170 ;
        RECT 1111.630 -9.260 1112.810 -8.080 ;
        RECT 1113.230 -9.260 1114.410 -8.080 ;
        RECT 1111.630 -10.860 1112.810 -9.680 ;
        RECT 1113.230 -10.860 1114.410 -9.680 ;
        RECT 1291.630 3529.360 1292.810 3530.540 ;
        RECT 1293.230 3529.360 1294.410 3530.540 ;
        RECT 1291.630 3527.760 1292.810 3528.940 ;
        RECT 1293.230 3527.760 1294.410 3528.940 ;
        RECT 1291.630 3458.590 1292.810 3459.770 ;
        RECT 1293.230 3458.590 1294.410 3459.770 ;
        RECT 1291.630 3456.990 1292.810 3458.170 ;
        RECT 1293.230 3456.990 1294.410 3458.170 ;
        RECT 1291.630 3278.590 1292.810 3279.770 ;
        RECT 1293.230 3278.590 1294.410 3279.770 ;
        RECT 1291.630 3276.990 1292.810 3278.170 ;
        RECT 1293.230 3276.990 1294.410 3278.170 ;
        RECT 1291.630 3098.590 1292.810 3099.770 ;
        RECT 1293.230 3098.590 1294.410 3099.770 ;
        RECT 1291.630 3096.990 1292.810 3098.170 ;
        RECT 1293.230 3096.990 1294.410 3098.170 ;
        RECT 1291.630 2918.590 1292.810 2919.770 ;
        RECT 1293.230 2918.590 1294.410 2919.770 ;
        RECT 1291.630 2916.990 1292.810 2918.170 ;
        RECT 1293.230 2916.990 1294.410 2918.170 ;
        RECT 1291.630 2738.590 1292.810 2739.770 ;
        RECT 1293.230 2738.590 1294.410 2739.770 ;
        RECT 1291.630 2736.990 1292.810 2738.170 ;
        RECT 1293.230 2736.990 1294.410 2738.170 ;
        RECT 1291.630 2558.590 1292.810 2559.770 ;
        RECT 1293.230 2558.590 1294.410 2559.770 ;
        RECT 1291.630 2556.990 1292.810 2558.170 ;
        RECT 1293.230 2556.990 1294.410 2558.170 ;
        RECT 1291.630 2378.590 1292.810 2379.770 ;
        RECT 1293.230 2378.590 1294.410 2379.770 ;
        RECT 1291.630 2376.990 1292.810 2378.170 ;
        RECT 1293.230 2376.990 1294.410 2378.170 ;
        RECT 1291.630 2198.590 1292.810 2199.770 ;
        RECT 1293.230 2198.590 1294.410 2199.770 ;
        RECT 1291.630 2196.990 1292.810 2198.170 ;
        RECT 1293.230 2196.990 1294.410 2198.170 ;
        RECT 1291.630 2018.590 1292.810 2019.770 ;
        RECT 1293.230 2018.590 1294.410 2019.770 ;
        RECT 1291.630 2016.990 1292.810 2018.170 ;
        RECT 1293.230 2016.990 1294.410 2018.170 ;
        RECT 1291.630 1838.590 1292.810 1839.770 ;
        RECT 1293.230 1838.590 1294.410 1839.770 ;
        RECT 1291.630 1836.990 1292.810 1838.170 ;
        RECT 1293.230 1836.990 1294.410 1838.170 ;
        RECT 1291.630 1658.590 1292.810 1659.770 ;
        RECT 1293.230 1658.590 1294.410 1659.770 ;
        RECT 1291.630 1656.990 1292.810 1658.170 ;
        RECT 1293.230 1656.990 1294.410 1658.170 ;
        RECT 1291.630 1478.590 1292.810 1479.770 ;
        RECT 1293.230 1478.590 1294.410 1479.770 ;
        RECT 1291.630 1476.990 1292.810 1478.170 ;
        RECT 1293.230 1476.990 1294.410 1478.170 ;
        RECT 1291.630 1298.590 1292.810 1299.770 ;
        RECT 1293.230 1298.590 1294.410 1299.770 ;
        RECT 1291.630 1296.990 1292.810 1298.170 ;
        RECT 1293.230 1296.990 1294.410 1298.170 ;
        RECT 1291.630 1118.590 1292.810 1119.770 ;
        RECT 1293.230 1118.590 1294.410 1119.770 ;
        RECT 1291.630 1116.990 1292.810 1118.170 ;
        RECT 1293.230 1116.990 1294.410 1118.170 ;
        RECT 1291.630 938.590 1292.810 939.770 ;
        RECT 1293.230 938.590 1294.410 939.770 ;
        RECT 1291.630 936.990 1292.810 938.170 ;
        RECT 1293.230 936.990 1294.410 938.170 ;
        RECT 1291.630 758.590 1292.810 759.770 ;
        RECT 1293.230 758.590 1294.410 759.770 ;
        RECT 1291.630 756.990 1292.810 758.170 ;
        RECT 1293.230 756.990 1294.410 758.170 ;
        RECT 1291.630 578.590 1292.810 579.770 ;
        RECT 1293.230 578.590 1294.410 579.770 ;
        RECT 1291.630 576.990 1292.810 578.170 ;
        RECT 1293.230 576.990 1294.410 578.170 ;
        RECT 1291.630 398.590 1292.810 399.770 ;
        RECT 1293.230 398.590 1294.410 399.770 ;
        RECT 1291.630 396.990 1292.810 398.170 ;
        RECT 1293.230 396.990 1294.410 398.170 ;
        RECT 1291.630 218.590 1292.810 219.770 ;
        RECT 1293.230 218.590 1294.410 219.770 ;
        RECT 1291.630 216.990 1292.810 218.170 ;
        RECT 1293.230 216.990 1294.410 218.170 ;
        RECT 1291.630 38.590 1292.810 39.770 ;
        RECT 1293.230 38.590 1294.410 39.770 ;
        RECT 1291.630 36.990 1292.810 38.170 ;
        RECT 1293.230 36.990 1294.410 38.170 ;
        RECT 1291.630 -9.260 1292.810 -8.080 ;
        RECT 1293.230 -9.260 1294.410 -8.080 ;
        RECT 1291.630 -10.860 1292.810 -9.680 ;
        RECT 1293.230 -10.860 1294.410 -9.680 ;
        RECT 1471.630 3529.360 1472.810 3530.540 ;
        RECT 1473.230 3529.360 1474.410 3530.540 ;
        RECT 1471.630 3527.760 1472.810 3528.940 ;
        RECT 1473.230 3527.760 1474.410 3528.940 ;
        RECT 1471.630 3458.590 1472.810 3459.770 ;
        RECT 1473.230 3458.590 1474.410 3459.770 ;
        RECT 1471.630 3456.990 1472.810 3458.170 ;
        RECT 1473.230 3456.990 1474.410 3458.170 ;
        RECT 1471.630 3278.590 1472.810 3279.770 ;
        RECT 1473.230 3278.590 1474.410 3279.770 ;
        RECT 1471.630 3276.990 1472.810 3278.170 ;
        RECT 1473.230 3276.990 1474.410 3278.170 ;
        RECT 1471.630 3098.590 1472.810 3099.770 ;
        RECT 1473.230 3098.590 1474.410 3099.770 ;
        RECT 1471.630 3096.990 1472.810 3098.170 ;
        RECT 1473.230 3096.990 1474.410 3098.170 ;
        RECT 1471.630 2918.590 1472.810 2919.770 ;
        RECT 1473.230 2918.590 1474.410 2919.770 ;
        RECT 1471.630 2916.990 1472.810 2918.170 ;
        RECT 1473.230 2916.990 1474.410 2918.170 ;
        RECT 1471.630 2738.590 1472.810 2739.770 ;
        RECT 1473.230 2738.590 1474.410 2739.770 ;
        RECT 1471.630 2736.990 1472.810 2738.170 ;
        RECT 1473.230 2736.990 1474.410 2738.170 ;
        RECT 1471.630 2558.590 1472.810 2559.770 ;
        RECT 1473.230 2558.590 1474.410 2559.770 ;
        RECT 1471.630 2556.990 1472.810 2558.170 ;
        RECT 1473.230 2556.990 1474.410 2558.170 ;
        RECT 1471.630 2378.590 1472.810 2379.770 ;
        RECT 1473.230 2378.590 1474.410 2379.770 ;
        RECT 1471.630 2376.990 1472.810 2378.170 ;
        RECT 1473.230 2376.990 1474.410 2378.170 ;
        RECT 1471.630 2198.590 1472.810 2199.770 ;
        RECT 1473.230 2198.590 1474.410 2199.770 ;
        RECT 1471.630 2196.990 1472.810 2198.170 ;
        RECT 1473.230 2196.990 1474.410 2198.170 ;
        RECT 1471.630 2018.590 1472.810 2019.770 ;
        RECT 1473.230 2018.590 1474.410 2019.770 ;
        RECT 1471.630 2016.990 1472.810 2018.170 ;
        RECT 1473.230 2016.990 1474.410 2018.170 ;
        RECT 1471.630 1838.590 1472.810 1839.770 ;
        RECT 1473.230 1838.590 1474.410 1839.770 ;
        RECT 1471.630 1836.990 1472.810 1838.170 ;
        RECT 1473.230 1836.990 1474.410 1838.170 ;
        RECT 1471.630 1658.590 1472.810 1659.770 ;
        RECT 1473.230 1658.590 1474.410 1659.770 ;
        RECT 1471.630 1656.990 1472.810 1658.170 ;
        RECT 1473.230 1656.990 1474.410 1658.170 ;
        RECT 1471.630 1478.590 1472.810 1479.770 ;
        RECT 1473.230 1478.590 1474.410 1479.770 ;
        RECT 1471.630 1476.990 1472.810 1478.170 ;
        RECT 1473.230 1476.990 1474.410 1478.170 ;
        RECT 1471.630 1298.590 1472.810 1299.770 ;
        RECT 1473.230 1298.590 1474.410 1299.770 ;
        RECT 1471.630 1296.990 1472.810 1298.170 ;
        RECT 1473.230 1296.990 1474.410 1298.170 ;
        RECT 1471.630 1118.590 1472.810 1119.770 ;
        RECT 1473.230 1118.590 1474.410 1119.770 ;
        RECT 1471.630 1116.990 1472.810 1118.170 ;
        RECT 1473.230 1116.990 1474.410 1118.170 ;
        RECT 1471.630 938.590 1472.810 939.770 ;
        RECT 1473.230 938.590 1474.410 939.770 ;
        RECT 1471.630 936.990 1472.810 938.170 ;
        RECT 1473.230 936.990 1474.410 938.170 ;
        RECT 1471.630 758.590 1472.810 759.770 ;
        RECT 1473.230 758.590 1474.410 759.770 ;
        RECT 1471.630 756.990 1472.810 758.170 ;
        RECT 1473.230 756.990 1474.410 758.170 ;
        RECT 1471.630 578.590 1472.810 579.770 ;
        RECT 1473.230 578.590 1474.410 579.770 ;
        RECT 1471.630 576.990 1472.810 578.170 ;
        RECT 1473.230 576.990 1474.410 578.170 ;
        RECT 1471.630 398.590 1472.810 399.770 ;
        RECT 1473.230 398.590 1474.410 399.770 ;
        RECT 1471.630 396.990 1472.810 398.170 ;
        RECT 1473.230 396.990 1474.410 398.170 ;
        RECT 1471.630 218.590 1472.810 219.770 ;
        RECT 1473.230 218.590 1474.410 219.770 ;
        RECT 1471.630 216.990 1472.810 218.170 ;
        RECT 1473.230 216.990 1474.410 218.170 ;
        RECT 1471.630 38.590 1472.810 39.770 ;
        RECT 1473.230 38.590 1474.410 39.770 ;
        RECT 1471.630 36.990 1472.810 38.170 ;
        RECT 1473.230 36.990 1474.410 38.170 ;
        RECT 1471.630 -9.260 1472.810 -8.080 ;
        RECT 1473.230 -9.260 1474.410 -8.080 ;
        RECT 1471.630 -10.860 1472.810 -9.680 ;
        RECT 1473.230 -10.860 1474.410 -9.680 ;
        RECT 1651.630 3529.360 1652.810 3530.540 ;
        RECT 1653.230 3529.360 1654.410 3530.540 ;
        RECT 1651.630 3527.760 1652.810 3528.940 ;
        RECT 1653.230 3527.760 1654.410 3528.940 ;
        RECT 1651.630 3458.590 1652.810 3459.770 ;
        RECT 1653.230 3458.590 1654.410 3459.770 ;
        RECT 1651.630 3456.990 1652.810 3458.170 ;
        RECT 1653.230 3456.990 1654.410 3458.170 ;
        RECT 1651.630 3278.590 1652.810 3279.770 ;
        RECT 1653.230 3278.590 1654.410 3279.770 ;
        RECT 1651.630 3276.990 1652.810 3278.170 ;
        RECT 1653.230 3276.990 1654.410 3278.170 ;
        RECT 1651.630 3098.590 1652.810 3099.770 ;
        RECT 1653.230 3098.590 1654.410 3099.770 ;
        RECT 1651.630 3096.990 1652.810 3098.170 ;
        RECT 1653.230 3096.990 1654.410 3098.170 ;
        RECT 1651.630 2918.590 1652.810 2919.770 ;
        RECT 1653.230 2918.590 1654.410 2919.770 ;
        RECT 1651.630 2916.990 1652.810 2918.170 ;
        RECT 1653.230 2916.990 1654.410 2918.170 ;
        RECT 1651.630 2738.590 1652.810 2739.770 ;
        RECT 1653.230 2738.590 1654.410 2739.770 ;
        RECT 1651.630 2736.990 1652.810 2738.170 ;
        RECT 1653.230 2736.990 1654.410 2738.170 ;
        RECT 1651.630 2558.590 1652.810 2559.770 ;
        RECT 1653.230 2558.590 1654.410 2559.770 ;
        RECT 1651.630 2556.990 1652.810 2558.170 ;
        RECT 1653.230 2556.990 1654.410 2558.170 ;
        RECT 1651.630 2378.590 1652.810 2379.770 ;
        RECT 1653.230 2378.590 1654.410 2379.770 ;
        RECT 1651.630 2376.990 1652.810 2378.170 ;
        RECT 1653.230 2376.990 1654.410 2378.170 ;
        RECT 1651.630 2198.590 1652.810 2199.770 ;
        RECT 1653.230 2198.590 1654.410 2199.770 ;
        RECT 1651.630 2196.990 1652.810 2198.170 ;
        RECT 1653.230 2196.990 1654.410 2198.170 ;
        RECT 1651.630 2018.590 1652.810 2019.770 ;
        RECT 1653.230 2018.590 1654.410 2019.770 ;
        RECT 1651.630 2016.990 1652.810 2018.170 ;
        RECT 1653.230 2016.990 1654.410 2018.170 ;
        RECT 1651.630 1838.590 1652.810 1839.770 ;
        RECT 1653.230 1838.590 1654.410 1839.770 ;
        RECT 1651.630 1836.990 1652.810 1838.170 ;
        RECT 1653.230 1836.990 1654.410 1838.170 ;
        RECT 1651.630 1658.590 1652.810 1659.770 ;
        RECT 1653.230 1658.590 1654.410 1659.770 ;
        RECT 1651.630 1656.990 1652.810 1658.170 ;
        RECT 1653.230 1656.990 1654.410 1658.170 ;
        RECT 1651.630 1478.590 1652.810 1479.770 ;
        RECT 1653.230 1478.590 1654.410 1479.770 ;
        RECT 1651.630 1476.990 1652.810 1478.170 ;
        RECT 1653.230 1476.990 1654.410 1478.170 ;
        RECT 1651.630 1298.590 1652.810 1299.770 ;
        RECT 1653.230 1298.590 1654.410 1299.770 ;
        RECT 1651.630 1296.990 1652.810 1298.170 ;
        RECT 1653.230 1296.990 1654.410 1298.170 ;
        RECT 1651.630 1118.590 1652.810 1119.770 ;
        RECT 1653.230 1118.590 1654.410 1119.770 ;
        RECT 1651.630 1116.990 1652.810 1118.170 ;
        RECT 1653.230 1116.990 1654.410 1118.170 ;
        RECT 1651.630 938.590 1652.810 939.770 ;
        RECT 1653.230 938.590 1654.410 939.770 ;
        RECT 1651.630 936.990 1652.810 938.170 ;
        RECT 1653.230 936.990 1654.410 938.170 ;
        RECT 1651.630 758.590 1652.810 759.770 ;
        RECT 1653.230 758.590 1654.410 759.770 ;
        RECT 1651.630 756.990 1652.810 758.170 ;
        RECT 1653.230 756.990 1654.410 758.170 ;
        RECT 1651.630 578.590 1652.810 579.770 ;
        RECT 1653.230 578.590 1654.410 579.770 ;
        RECT 1651.630 576.990 1652.810 578.170 ;
        RECT 1653.230 576.990 1654.410 578.170 ;
        RECT 1651.630 398.590 1652.810 399.770 ;
        RECT 1653.230 398.590 1654.410 399.770 ;
        RECT 1651.630 396.990 1652.810 398.170 ;
        RECT 1653.230 396.990 1654.410 398.170 ;
        RECT 1651.630 218.590 1652.810 219.770 ;
        RECT 1653.230 218.590 1654.410 219.770 ;
        RECT 1651.630 216.990 1652.810 218.170 ;
        RECT 1653.230 216.990 1654.410 218.170 ;
        RECT 1651.630 38.590 1652.810 39.770 ;
        RECT 1653.230 38.590 1654.410 39.770 ;
        RECT 1651.630 36.990 1652.810 38.170 ;
        RECT 1653.230 36.990 1654.410 38.170 ;
        RECT 1651.630 -9.260 1652.810 -8.080 ;
        RECT 1653.230 -9.260 1654.410 -8.080 ;
        RECT 1651.630 -10.860 1652.810 -9.680 ;
        RECT 1653.230 -10.860 1654.410 -9.680 ;
        RECT 1831.630 3529.360 1832.810 3530.540 ;
        RECT 1833.230 3529.360 1834.410 3530.540 ;
        RECT 1831.630 3527.760 1832.810 3528.940 ;
        RECT 1833.230 3527.760 1834.410 3528.940 ;
        RECT 1831.630 3458.590 1832.810 3459.770 ;
        RECT 1833.230 3458.590 1834.410 3459.770 ;
        RECT 1831.630 3456.990 1832.810 3458.170 ;
        RECT 1833.230 3456.990 1834.410 3458.170 ;
        RECT 1831.630 3278.590 1832.810 3279.770 ;
        RECT 1833.230 3278.590 1834.410 3279.770 ;
        RECT 1831.630 3276.990 1832.810 3278.170 ;
        RECT 1833.230 3276.990 1834.410 3278.170 ;
        RECT 1831.630 3098.590 1832.810 3099.770 ;
        RECT 1833.230 3098.590 1834.410 3099.770 ;
        RECT 1831.630 3096.990 1832.810 3098.170 ;
        RECT 1833.230 3096.990 1834.410 3098.170 ;
        RECT 1831.630 2918.590 1832.810 2919.770 ;
        RECT 1833.230 2918.590 1834.410 2919.770 ;
        RECT 1831.630 2916.990 1832.810 2918.170 ;
        RECT 1833.230 2916.990 1834.410 2918.170 ;
        RECT 1831.630 2738.590 1832.810 2739.770 ;
        RECT 1833.230 2738.590 1834.410 2739.770 ;
        RECT 1831.630 2736.990 1832.810 2738.170 ;
        RECT 1833.230 2736.990 1834.410 2738.170 ;
        RECT 1831.630 2558.590 1832.810 2559.770 ;
        RECT 1833.230 2558.590 1834.410 2559.770 ;
        RECT 1831.630 2556.990 1832.810 2558.170 ;
        RECT 1833.230 2556.990 1834.410 2558.170 ;
        RECT 1831.630 2378.590 1832.810 2379.770 ;
        RECT 1833.230 2378.590 1834.410 2379.770 ;
        RECT 1831.630 2376.990 1832.810 2378.170 ;
        RECT 1833.230 2376.990 1834.410 2378.170 ;
        RECT 1831.630 2198.590 1832.810 2199.770 ;
        RECT 1833.230 2198.590 1834.410 2199.770 ;
        RECT 1831.630 2196.990 1832.810 2198.170 ;
        RECT 1833.230 2196.990 1834.410 2198.170 ;
        RECT 1831.630 2018.590 1832.810 2019.770 ;
        RECT 1833.230 2018.590 1834.410 2019.770 ;
        RECT 1831.630 2016.990 1832.810 2018.170 ;
        RECT 1833.230 2016.990 1834.410 2018.170 ;
        RECT 1831.630 1838.590 1832.810 1839.770 ;
        RECT 1833.230 1838.590 1834.410 1839.770 ;
        RECT 1831.630 1836.990 1832.810 1838.170 ;
        RECT 1833.230 1836.990 1834.410 1838.170 ;
        RECT 1831.630 1658.590 1832.810 1659.770 ;
        RECT 1833.230 1658.590 1834.410 1659.770 ;
        RECT 1831.630 1656.990 1832.810 1658.170 ;
        RECT 1833.230 1656.990 1834.410 1658.170 ;
        RECT 1831.630 1478.590 1832.810 1479.770 ;
        RECT 1833.230 1478.590 1834.410 1479.770 ;
        RECT 1831.630 1476.990 1832.810 1478.170 ;
        RECT 1833.230 1476.990 1834.410 1478.170 ;
        RECT 1831.630 1298.590 1832.810 1299.770 ;
        RECT 1833.230 1298.590 1834.410 1299.770 ;
        RECT 1831.630 1296.990 1832.810 1298.170 ;
        RECT 1833.230 1296.990 1834.410 1298.170 ;
        RECT 1831.630 1118.590 1832.810 1119.770 ;
        RECT 1833.230 1118.590 1834.410 1119.770 ;
        RECT 1831.630 1116.990 1832.810 1118.170 ;
        RECT 1833.230 1116.990 1834.410 1118.170 ;
        RECT 1831.630 938.590 1832.810 939.770 ;
        RECT 1833.230 938.590 1834.410 939.770 ;
        RECT 1831.630 936.990 1832.810 938.170 ;
        RECT 1833.230 936.990 1834.410 938.170 ;
        RECT 1831.630 758.590 1832.810 759.770 ;
        RECT 1833.230 758.590 1834.410 759.770 ;
        RECT 1831.630 756.990 1832.810 758.170 ;
        RECT 1833.230 756.990 1834.410 758.170 ;
        RECT 1831.630 578.590 1832.810 579.770 ;
        RECT 1833.230 578.590 1834.410 579.770 ;
        RECT 1831.630 576.990 1832.810 578.170 ;
        RECT 1833.230 576.990 1834.410 578.170 ;
        RECT 1831.630 398.590 1832.810 399.770 ;
        RECT 1833.230 398.590 1834.410 399.770 ;
        RECT 1831.630 396.990 1832.810 398.170 ;
        RECT 1833.230 396.990 1834.410 398.170 ;
        RECT 1831.630 218.590 1832.810 219.770 ;
        RECT 1833.230 218.590 1834.410 219.770 ;
        RECT 1831.630 216.990 1832.810 218.170 ;
        RECT 1833.230 216.990 1834.410 218.170 ;
        RECT 1831.630 38.590 1832.810 39.770 ;
        RECT 1833.230 38.590 1834.410 39.770 ;
        RECT 1831.630 36.990 1832.810 38.170 ;
        RECT 1833.230 36.990 1834.410 38.170 ;
        RECT 1831.630 -9.260 1832.810 -8.080 ;
        RECT 1833.230 -9.260 1834.410 -8.080 ;
        RECT 1831.630 -10.860 1832.810 -9.680 ;
        RECT 1833.230 -10.860 1834.410 -9.680 ;
        RECT 2011.630 3529.360 2012.810 3530.540 ;
        RECT 2013.230 3529.360 2014.410 3530.540 ;
        RECT 2011.630 3527.760 2012.810 3528.940 ;
        RECT 2013.230 3527.760 2014.410 3528.940 ;
        RECT 2011.630 3458.590 2012.810 3459.770 ;
        RECT 2013.230 3458.590 2014.410 3459.770 ;
        RECT 2011.630 3456.990 2012.810 3458.170 ;
        RECT 2013.230 3456.990 2014.410 3458.170 ;
        RECT 2011.630 3278.590 2012.810 3279.770 ;
        RECT 2013.230 3278.590 2014.410 3279.770 ;
        RECT 2011.630 3276.990 2012.810 3278.170 ;
        RECT 2013.230 3276.990 2014.410 3278.170 ;
        RECT 2011.630 3098.590 2012.810 3099.770 ;
        RECT 2013.230 3098.590 2014.410 3099.770 ;
        RECT 2011.630 3096.990 2012.810 3098.170 ;
        RECT 2013.230 3096.990 2014.410 3098.170 ;
        RECT 2011.630 2918.590 2012.810 2919.770 ;
        RECT 2013.230 2918.590 2014.410 2919.770 ;
        RECT 2011.630 2916.990 2012.810 2918.170 ;
        RECT 2013.230 2916.990 2014.410 2918.170 ;
        RECT 2011.630 2738.590 2012.810 2739.770 ;
        RECT 2013.230 2738.590 2014.410 2739.770 ;
        RECT 2011.630 2736.990 2012.810 2738.170 ;
        RECT 2013.230 2736.990 2014.410 2738.170 ;
        RECT 2011.630 2558.590 2012.810 2559.770 ;
        RECT 2013.230 2558.590 2014.410 2559.770 ;
        RECT 2011.630 2556.990 2012.810 2558.170 ;
        RECT 2013.230 2556.990 2014.410 2558.170 ;
        RECT 2011.630 2378.590 2012.810 2379.770 ;
        RECT 2013.230 2378.590 2014.410 2379.770 ;
        RECT 2011.630 2376.990 2012.810 2378.170 ;
        RECT 2013.230 2376.990 2014.410 2378.170 ;
        RECT 2011.630 2198.590 2012.810 2199.770 ;
        RECT 2013.230 2198.590 2014.410 2199.770 ;
        RECT 2011.630 2196.990 2012.810 2198.170 ;
        RECT 2013.230 2196.990 2014.410 2198.170 ;
        RECT 2011.630 2018.590 2012.810 2019.770 ;
        RECT 2013.230 2018.590 2014.410 2019.770 ;
        RECT 2011.630 2016.990 2012.810 2018.170 ;
        RECT 2013.230 2016.990 2014.410 2018.170 ;
        RECT 2011.630 1838.590 2012.810 1839.770 ;
        RECT 2013.230 1838.590 2014.410 1839.770 ;
        RECT 2011.630 1836.990 2012.810 1838.170 ;
        RECT 2013.230 1836.990 2014.410 1838.170 ;
        RECT 2011.630 1658.590 2012.810 1659.770 ;
        RECT 2013.230 1658.590 2014.410 1659.770 ;
        RECT 2011.630 1656.990 2012.810 1658.170 ;
        RECT 2013.230 1656.990 2014.410 1658.170 ;
        RECT 2011.630 1478.590 2012.810 1479.770 ;
        RECT 2013.230 1478.590 2014.410 1479.770 ;
        RECT 2011.630 1476.990 2012.810 1478.170 ;
        RECT 2013.230 1476.990 2014.410 1478.170 ;
        RECT 2011.630 1298.590 2012.810 1299.770 ;
        RECT 2013.230 1298.590 2014.410 1299.770 ;
        RECT 2011.630 1296.990 2012.810 1298.170 ;
        RECT 2013.230 1296.990 2014.410 1298.170 ;
        RECT 2011.630 1118.590 2012.810 1119.770 ;
        RECT 2013.230 1118.590 2014.410 1119.770 ;
        RECT 2011.630 1116.990 2012.810 1118.170 ;
        RECT 2013.230 1116.990 2014.410 1118.170 ;
        RECT 2011.630 938.590 2012.810 939.770 ;
        RECT 2013.230 938.590 2014.410 939.770 ;
        RECT 2011.630 936.990 2012.810 938.170 ;
        RECT 2013.230 936.990 2014.410 938.170 ;
        RECT 2011.630 758.590 2012.810 759.770 ;
        RECT 2013.230 758.590 2014.410 759.770 ;
        RECT 2011.630 756.990 2012.810 758.170 ;
        RECT 2013.230 756.990 2014.410 758.170 ;
        RECT 2011.630 578.590 2012.810 579.770 ;
        RECT 2013.230 578.590 2014.410 579.770 ;
        RECT 2011.630 576.990 2012.810 578.170 ;
        RECT 2013.230 576.990 2014.410 578.170 ;
        RECT 2011.630 398.590 2012.810 399.770 ;
        RECT 2013.230 398.590 2014.410 399.770 ;
        RECT 2011.630 396.990 2012.810 398.170 ;
        RECT 2013.230 396.990 2014.410 398.170 ;
        RECT 2011.630 218.590 2012.810 219.770 ;
        RECT 2013.230 218.590 2014.410 219.770 ;
        RECT 2011.630 216.990 2012.810 218.170 ;
        RECT 2013.230 216.990 2014.410 218.170 ;
        RECT 2011.630 38.590 2012.810 39.770 ;
        RECT 2013.230 38.590 2014.410 39.770 ;
        RECT 2011.630 36.990 2012.810 38.170 ;
        RECT 2013.230 36.990 2014.410 38.170 ;
        RECT 2011.630 -9.260 2012.810 -8.080 ;
        RECT 2013.230 -9.260 2014.410 -8.080 ;
        RECT 2011.630 -10.860 2012.810 -9.680 ;
        RECT 2013.230 -10.860 2014.410 -9.680 ;
        RECT 2191.630 3529.360 2192.810 3530.540 ;
        RECT 2193.230 3529.360 2194.410 3530.540 ;
        RECT 2191.630 3527.760 2192.810 3528.940 ;
        RECT 2193.230 3527.760 2194.410 3528.940 ;
        RECT 2191.630 3458.590 2192.810 3459.770 ;
        RECT 2193.230 3458.590 2194.410 3459.770 ;
        RECT 2191.630 3456.990 2192.810 3458.170 ;
        RECT 2193.230 3456.990 2194.410 3458.170 ;
        RECT 2191.630 3278.590 2192.810 3279.770 ;
        RECT 2193.230 3278.590 2194.410 3279.770 ;
        RECT 2191.630 3276.990 2192.810 3278.170 ;
        RECT 2193.230 3276.990 2194.410 3278.170 ;
        RECT 2191.630 3098.590 2192.810 3099.770 ;
        RECT 2193.230 3098.590 2194.410 3099.770 ;
        RECT 2191.630 3096.990 2192.810 3098.170 ;
        RECT 2193.230 3096.990 2194.410 3098.170 ;
        RECT 2191.630 2918.590 2192.810 2919.770 ;
        RECT 2193.230 2918.590 2194.410 2919.770 ;
        RECT 2191.630 2916.990 2192.810 2918.170 ;
        RECT 2193.230 2916.990 2194.410 2918.170 ;
        RECT 2191.630 2738.590 2192.810 2739.770 ;
        RECT 2193.230 2738.590 2194.410 2739.770 ;
        RECT 2191.630 2736.990 2192.810 2738.170 ;
        RECT 2193.230 2736.990 2194.410 2738.170 ;
        RECT 2191.630 2558.590 2192.810 2559.770 ;
        RECT 2193.230 2558.590 2194.410 2559.770 ;
        RECT 2191.630 2556.990 2192.810 2558.170 ;
        RECT 2193.230 2556.990 2194.410 2558.170 ;
        RECT 2191.630 2378.590 2192.810 2379.770 ;
        RECT 2193.230 2378.590 2194.410 2379.770 ;
        RECT 2191.630 2376.990 2192.810 2378.170 ;
        RECT 2193.230 2376.990 2194.410 2378.170 ;
        RECT 2191.630 2198.590 2192.810 2199.770 ;
        RECT 2193.230 2198.590 2194.410 2199.770 ;
        RECT 2191.630 2196.990 2192.810 2198.170 ;
        RECT 2193.230 2196.990 2194.410 2198.170 ;
        RECT 2191.630 2018.590 2192.810 2019.770 ;
        RECT 2193.230 2018.590 2194.410 2019.770 ;
        RECT 2191.630 2016.990 2192.810 2018.170 ;
        RECT 2193.230 2016.990 2194.410 2018.170 ;
        RECT 2191.630 1838.590 2192.810 1839.770 ;
        RECT 2193.230 1838.590 2194.410 1839.770 ;
        RECT 2191.630 1836.990 2192.810 1838.170 ;
        RECT 2193.230 1836.990 2194.410 1838.170 ;
        RECT 2191.630 1658.590 2192.810 1659.770 ;
        RECT 2193.230 1658.590 2194.410 1659.770 ;
        RECT 2191.630 1656.990 2192.810 1658.170 ;
        RECT 2193.230 1656.990 2194.410 1658.170 ;
        RECT 2191.630 1478.590 2192.810 1479.770 ;
        RECT 2193.230 1478.590 2194.410 1479.770 ;
        RECT 2191.630 1476.990 2192.810 1478.170 ;
        RECT 2193.230 1476.990 2194.410 1478.170 ;
        RECT 2191.630 1298.590 2192.810 1299.770 ;
        RECT 2193.230 1298.590 2194.410 1299.770 ;
        RECT 2191.630 1296.990 2192.810 1298.170 ;
        RECT 2193.230 1296.990 2194.410 1298.170 ;
        RECT 2191.630 1118.590 2192.810 1119.770 ;
        RECT 2193.230 1118.590 2194.410 1119.770 ;
        RECT 2191.630 1116.990 2192.810 1118.170 ;
        RECT 2193.230 1116.990 2194.410 1118.170 ;
        RECT 2191.630 938.590 2192.810 939.770 ;
        RECT 2193.230 938.590 2194.410 939.770 ;
        RECT 2191.630 936.990 2192.810 938.170 ;
        RECT 2193.230 936.990 2194.410 938.170 ;
        RECT 2191.630 758.590 2192.810 759.770 ;
        RECT 2193.230 758.590 2194.410 759.770 ;
        RECT 2191.630 756.990 2192.810 758.170 ;
        RECT 2193.230 756.990 2194.410 758.170 ;
        RECT 2191.630 578.590 2192.810 579.770 ;
        RECT 2193.230 578.590 2194.410 579.770 ;
        RECT 2191.630 576.990 2192.810 578.170 ;
        RECT 2193.230 576.990 2194.410 578.170 ;
        RECT 2191.630 398.590 2192.810 399.770 ;
        RECT 2193.230 398.590 2194.410 399.770 ;
        RECT 2191.630 396.990 2192.810 398.170 ;
        RECT 2193.230 396.990 2194.410 398.170 ;
        RECT 2191.630 218.590 2192.810 219.770 ;
        RECT 2193.230 218.590 2194.410 219.770 ;
        RECT 2191.630 216.990 2192.810 218.170 ;
        RECT 2193.230 216.990 2194.410 218.170 ;
        RECT 2191.630 38.590 2192.810 39.770 ;
        RECT 2193.230 38.590 2194.410 39.770 ;
        RECT 2191.630 36.990 2192.810 38.170 ;
        RECT 2193.230 36.990 2194.410 38.170 ;
        RECT 2191.630 -9.260 2192.810 -8.080 ;
        RECT 2193.230 -9.260 2194.410 -8.080 ;
        RECT 2191.630 -10.860 2192.810 -9.680 ;
        RECT 2193.230 -10.860 2194.410 -9.680 ;
        RECT 2371.630 3529.360 2372.810 3530.540 ;
        RECT 2373.230 3529.360 2374.410 3530.540 ;
        RECT 2371.630 3527.760 2372.810 3528.940 ;
        RECT 2373.230 3527.760 2374.410 3528.940 ;
        RECT 2371.630 3458.590 2372.810 3459.770 ;
        RECT 2373.230 3458.590 2374.410 3459.770 ;
        RECT 2371.630 3456.990 2372.810 3458.170 ;
        RECT 2373.230 3456.990 2374.410 3458.170 ;
        RECT 2371.630 3278.590 2372.810 3279.770 ;
        RECT 2373.230 3278.590 2374.410 3279.770 ;
        RECT 2371.630 3276.990 2372.810 3278.170 ;
        RECT 2373.230 3276.990 2374.410 3278.170 ;
        RECT 2371.630 3098.590 2372.810 3099.770 ;
        RECT 2373.230 3098.590 2374.410 3099.770 ;
        RECT 2371.630 3096.990 2372.810 3098.170 ;
        RECT 2373.230 3096.990 2374.410 3098.170 ;
        RECT 2371.630 2918.590 2372.810 2919.770 ;
        RECT 2373.230 2918.590 2374.410 2919.770 ;
        RECT 2371.630 2916.990 2372.810 2918.170 ;
        RECT 2373.230 2916.990 2374.410 2918.170 ;
        RECT 2371.630 2738.590 2372.810 2739.770 ;
        RECT 2373.230 2738.590 2374.410 2739.770 ;
        RECT 2371.630 2736.990 2372.810 2738.170 ;
        RECT 2373.230 2736.990 2374.410 2738.170 ;
        RECT 2371.630 2558.590 2372.810 2559.770 ;
        RECT 2373.230 2558.590 2374.410 2559.770 ;
        RECT 2371.630 2556.990 2372.810 2558.170 ;
        RECT 2373.230 2556.990 2374.410 2558.170 ;
        RECT 2371.630 2378.590 2372.810 2379.770 ;
        RECT 2373.230 2378.590 2374.410 2379.770 ;
        RECT 2371.630 2376.990 2372.810 2378.170 ;
        RECT 2373.230 2376.990 2374.410 2378.170 ;
        RECT 2371.630 2198.590 2372.810 2199.770 ;
        RECT 2373.230 2198.590 2374.410 2199.770 ;
        RECT 2371.630 2196.990 2372.810 2198.170 ;
        RECT 2373.230 2196.990 2374.410 2198.170 ;
        RECT 2371.630 2018.590 2372.810 2019.770 ;
        RECT 2373.230 2018.590 2374.410 2019.770 ;
        RECT 2371.630 2016.990 2372.810 2018.170 ;
        RECT 2373.230 2016.990 2374.410 2018.170 ;
        RECT 2371.630 1838.590 2372.810 1839.770 ;
        RECT 2373.230 1838.590 2374.410 1839.770 ;
        RECT 2371.630 1836.990 2372.810 1838.170 ;
        RECT 2373.230 1836.990 2374.410 1838.170 ;
        RECT 2371.630 1658.590 2372.810 1659.770 ;
        RECT 2373.230 1658.590 2374.410 1659.770 ;
        RECT 2371.630 1656.990 2372.810 1658.170 ;
        RECT 2373.230 1656.990 2374.410 1658.170 ;
        RECT 2371.630 1478.590 2372.810 1479.770 ;
        RECT 2373.230 1478.590 2374.410 1479.770 ;
        RECT 2371.630 1476.990 2372.810 1478.170 ;
        RECT 2373.230 1476.990 2374.410 1478.170 ;
        RECT 2371.630 1298.590 2372.810 1299.770 ;
        RECT 2373.230 1298.590 2374.410 1299.770 ;
        RECT 2371.630 1296.990 2372.810 1298.170 ;
        RECT 2373.230 1296.990 2374.410 1298.170 ;
        RECT 2371.630 1118.590 2372.810 1119.770 ;
        RECT 2373.230 1118.590 2374.410 1119.770 ;
        RECT 2371.630 1116.990 2372.810 1118.170 ;
        RECT 2373.230 1116.990 2374.410 1118.170 ;
        RECT 2371.630 938.590 2372.810 939.770 ;
        RECT 2373.230 938.590 2374.410 939.770 ;
        RECT 2371.630 936.990 2372.810 938.170 ;
        RECT 2373.230 936.990 2374.410 938.170 ;
        RECT 2371.630 758.590 2372.810 759.770 ;
        RECT 2373.230 758.590 2374.410 759.770 ;
        RECT 2371.630 756.990 2372.810 758.170 ;
        RECT 2373.230 756.990 2374.410 758.170 ;
        RECT 2371.630 578.590 2372.810 579.770 ;
        RECT 2373.230 578.590 2374.410 579.770 ;
        RECT 2371.630 576.990 2372.810 578.170 ;
        RECT 2373.230 576.990 2374.410 578.170 ;
        RECT 2371.630 398.590 2372.810 399.770 ;
        RECT 2373.230 398.590 2374.410 399.770 ;
        RECT 2371.630 396.990 2372.810 398.170 ;
        RECT 2373.230 396.990 2374.410 398.170 ;
        RECT 2371.630 218.590 2372.810 219.770 ;
        RECT 2373.230 218.590 2374.410 219.770 ;
        RECT 2371.630 216.990 2372.810 218.170 ;
        RECT 2373.230 216.990 2374.410 218.170 ;
        RECT 2371.630 38.590 2372.810 39.770 ;
        RECT 2373.230 38.590 2374.410 39.770 ;
        RECT 2371.630 36.990 2372.810 38.170 ;
        RECT 2373.230 36.990 2374.410 38.170 ;
        RECT 2371.630 -9.260 2372.810 -8.080 ;
        RECT 2373.230 -9.260 2374.410 -8.080 ;
        RECT 2371.630 -10.860 2372.810 -9.680 ;
        RECT 2373.230 -10.860 2374.410 -9.680 ;
        RECT 2551.630 3529.360 2552.810 3530.540 ;
        RECT 2553.230 3529.360 2554.410 3530.540 ;
        RECT 2551.630 3527.760 2552.810 3528.940 ;
        RECT 2553.230 3527.760 2554.410 3528.940 ;
        RECT 2551.630 3458.590 2552.810 3459.770 ;
        RECT 2553.230 3458.590 2554.410 3459.770 ;
        RECT 2551.630 3456.990 2552.810 3458.170 ;
        RECT 2553.230 3456.990 2554.410 3458.170 ;
        RECT 2551.630 3278.590 2552.810 3279.770 ;
        RECT 2553.230 3278.590 2554.410 3279.770 ;
        RECT 2551.630 3276.990 2552.810 3278.170 ;
        RECT 2553.230 3276.990 2554.410 3278.170 ;
        RECT 2551.630 3098.590 2552.810 3099.770 ;
        RECT 2553.230 3098.590 2554.410 3099.770 ;
        RECT 2551.630 3096.990 2552.810 3098.170 ;
        RECT 2553.230 3096.990 2554.410 3098.170 ;
        RECT 2551.630 2918.590 2552.810 2919.770 ;
        RECT 2553.230 2918.590 2554.410 2919.770 ;
        RECT 2551.630 2916.990 2552.810 2918.170 ;
        RECT 2553.230 2916.990 2554.410 2918.170 ;
        RECT 2551.630 2738.590 2552.810 2739.770 ;
        RECT 2553.230 2738.590 2554.410 2739.770 ;
        RECT 2551.630 2736.990 2552.810 2738.170 ;
        RECT 2553.230 2736.990 2554.410 2738.170 ;
        RECT 2551.630 2558.590 2552.810 2559.770 ;
        RECT 2553.230 2558.590 2554.410 2559.770 ;
        RECT 2551.630 2556.990 2552.810 2558.170 ;
        RECT 2553.230 2556.990 2554.410 2558.170 ;
        RECT 2551.630 2378.590 2552.810 2379.770 ;
        RECT 2553.230 2378.590 2554.410 2379.770 ;
        RECT 2551.630 2376.990 2552.810 2378.170 ;
        RECT 2553.230 2376.990 2554.410 2378.170 ;
        RECT 2551.630 2198.590 2552.810 2199.770 ;
        RECT 2553.230 2198.590 2554.410 2199.770 ;
        RECT 2551.630 2196.990 2552.810 2198.170 ;
        RECT 2553.230 2196.990 2554.410 2198.170 ;
        RECT 2551.630 2018.590 2552.810 2019.770 ;
        RECT 2553.230 2018.590 2554.410 2019.770 ;
        RECT 2551.630 2016.990 2552.810 2018.170 ;
        RECT 2553.230 2016.990 2554.410 2018.170 ;
        RECT 2551.630 1838.590 2552.810 1839.770 ;
        RECT 2553.230 1838.590 2554.410 1839.770 ;
        RECT 2551.630 1836.990 2552.810 1838.170 ;
        RECT 2553.230 1836.990 2554.410 1838.170 ;
        RECT 2551.630 1658.590 2552.810 1659.770 ;
        RECT 2553.230 1658.590 2554.410 1659.770 ;
        RECT 2551.630 1656.990 2552.810 1658.170 ;
        RECT 2553.230 1656.990 2554.410 1658.170 ;
        RECT 2551.630 1478.590 2552.810 1479.770 ;
        RECT 2553.230 1478.590 2554.410 1479.770 ;
        RECT 2551.630 1476.990 2552.810 1478.170 ;
        RECT 2553.230 1476.990 2554.410 1478.170 ;
        RECT 2551.630 1298.590 2552.810 1299.770 ;
        RECT 2553.230 1298.590 2554.410 1299.770 ;
        RECT 2551.630 1296.990 2552.810 1298.170 ;
        RECT 2553.230 1296.990 2554.410 1298.170 ;
        RECT 2551.630 1118.590 2552.810 1119.770 ;
        RECT 2553.230 1118.590 2554.410 1119.770 ;
        RECT 2551.630 1116.990 2552.810 1118.170 ;
        RECT 2553.230 1116.990 2554.410 1118.170 ;
        RECT 2551.630 938.590 2552.810 939.770 ;
        RECT 2553.230 938.590 2554.410 939.770 ;
        RECT 2551.630 936.990 2552.810 938.170 ;
        RECT 2553.230 936.990 2554.410 938.170 ;
        RECT 2551.630 758.590 2552.810 759.770 ;
        RECT 2553.230 758.590 2554.410 759.770 ;
        RECT 2551.630 756.990 2552.810 758.170 ;
        RECT 2553.230 756.990 2554.410 758.170 ;
        RECT 2551.630 578.590 2552.810 579.770 ;
        RECT 2553.230 578.590 2554.410 579.770 ;
        RECT 2551.630 576.990 2552.810 578.170 ;
        RECT 2553.230 576.990 2554.410 578.170 ;
        RECT 2551.630 398.590 2552.810 399.770 ;
        RECT 2553.230 398.590 2554.410 399.770 ;
        RECT 2551.630 396.990 2552.810 398.170 ;
        RECT 2553.230 396.990 2554.410 398.170 ;
        RECT 2551.630 218.590 2552.810 219.770 ;
        RECT 2553.230 218.590 2554.410 219.770 ;
        RECT 2551.630 216.990 2552.810 218.170 ;
        RECT 2553.230 216.990 2554.410 218.170 ;
        RECT 2551.630 38.590 2552.810 39.770 ;
        RECT 2553.230 38.590 2554.410 39.770 ;
        RECT 2551.630 36.990 2552.810 38.170 ;
        RECT 2553.230 36.990 2554.410 38.170 ;
        RECT 2551.630 -9.260 2552.810 -8.080 ;
        RECT 2553.230 -9.260 2554.410 -8.080 ;
        RECT 2551.630 -10.860 2552.810 -9.680 ;
        RECT 2553.230 -10.860 2554.410 -9.680 ;
        RECT 2731.630 3529.360 2732.810 3530.540 ;
        RECT 2733.230 3529.360 2734.410 3530.540 ;
        RECT 2731.630 3527.760 2732.810 3528.940 ;
        RECT 2733.230 3527.760 2734.410 3528.940 ;
        RECT 2731.630 3458.590 2732.810 3459.770 ;
        RECT 2733.230 3458.590 2734.410 3459.770 ;
        RECT 2731.630 3456.990 2732.810 3458.170 ;
        RECT 2733.230 3456.990 2734.410 3458.170 ;
        RECT 2731.630 3278.590 2732.810 3279.770 ;
        RECT 2733.230 3278.590 2734.410 3279.770 ;
        RECT 2731.630 3276.990 2732.810 3278.170 ;
        RECT 2733.230 3276.990 2734.410 3278.170 ;
        RECT 2731.630 3098.590 2732.810 3099.770 ;
        RECT 2733.230 3098.590 2734.410 3099.770 ;
        RECT 2731.630 3096.990 2732.810 3098.170 ;
        RECT 2733.230 3096.990 2734.410 3098.170 ;
        RECT 2731.630 2918.590 2732.810 2919.770 ;
        RECT 2733.230 2918.590 2734.410 2919.770 ;
        RECT 2731.630 2916.990 2732.810 2918.170 ;
        RECT 2733.230 2916.990 2734.410 2918.170 ;
        RECT 2731.630 2738.590 2732.810 2739.770 ;
        RECT 2733.230 2738.590 2734.410 2739.770 ;
        RECT 2731.630 2736.990 2732.810 2738.170 ;
        RECT 2733.230 2736.990 2734.410 2738.170 ;
        RECT 2731.630 2558.590 2732.810 2559.770 ;
        RECT 2733.230 2558.590 2734.410 2559.770 ;
        RECT 2731.630 2556.990 2732.810 2558.170 ;
        RECT 2733.230 2556.990 2734.410 2558.170 ;
        RECT 2731.630 2378.590 2732.810 2379.770 ;
        RECT 2733.230 2378.590 2734.410 2379.770 ;
        RECT 2731.630 2376.990 2732.810 2378.170 ;
        RECT 2733.230 2376.990 2734.410 2378.170 ;
        RECT 2731.630 2198.590 2732.810 2199.770 ;
        RECT 2733.230 2198.590 2734.410 2199.770 ;
        RECT 2731.630 2196.990 2732.810 2198.170 ;
        RECT 2733.230 2196.990 2734.410 2198.170 ;
        RECT 2731.630 2018.590 2732.810 2019.770 ;
        RECT 2733.230 2018.590 2734.410 2019.770 ;
        RECT 2731.630 2016.990 2732.810 2018.170 ;
        RECT 2733.230 2016.990 2734.410 2018.170 ;
        RECT 2731.630 1838.590 2732.810 1839.770 ;
        RECT 2733.230 1838.590 2734.410 1839.770 ;
        RECT 2731.630 1836.990 2732.810 1838.170 ;
        RECT 2733.230 1836.990 2734.410 1838.170 ;
        RECT 2731.630 1658.590 2732.810 1659.770 ;
        RECT 2733.230 1658.590 2734.410 1659.770 ;
        RECT 2731.630 1656.990 2732.810 1658.170 ;
        RECT 2733.230 1656.990 2734.410 1658.170 ;
        RECT 2731.630 1478.590 2732.810 1479.770 ;
        RECT 2733.230 1478.590 2734.410 1479.770 ;
        RECT 2731.630 1476.990 2732.810 1478.170 ;
        RECT 2733.230 1476.990 2734.410 1478.170 ;
        RECT 2731.630 1298.590 2732.810 1299.770 ;
        RECT 2733.230 1298.590 2734.410 1299.770 ;
        RECT 2731.630 1296.990 2732.810 1298.170 ;
        RECT 2733.230 1296.990 2734.410 1298.170 ;
        RECT 2731.630 1118.590 2732.810 1119.770 ;
        RECT 2733.230 1118.590 2734.410 1119.770 ;
        RECT 2731.630 1116.990 2732.810 1118.170 ;
        RECT 2733.230 1116.990 2734.410 1118.170 ;
        RECT 2731.630 938.590 2732.810 939.770 ;
        RECT 2733.230 938.590 2734.410 939.770 ;
        RECT 2731.630 936.990 2732.810 938.170 ;
        RECT 2733.230 936.990 2734.410 938.170 ;
        RECT 2731.630 758.590 2732.810 759.770 ;
        RECT 2733.230 758.590 2734.410 759.770 ;
        RECT 2731.630 756.990 2732.810 758.170 ;
        RECT 2733.230 756.990 2734.410 758.170 ;
        RECT 2731.630 578.590 2732.810 579.770 ;
        RECT 2733.230 578.590 2734.410 579.770 ;
        RECT 2731.630 576.990 2732.810 578.170 ;
        RECT 2733.230 576.990 2734.410 578.170 ;
        RECT 2731.630 398.590 2732.810 399.770 ;
        RECT 2733.230 398.590 2734.410 399.770 ;
        RECT 2731.630 396.990 2732.810 398.170 ;
        RECT 2733.230 396.990 2734.410 398.170 ;
        RECT 2731.630 218.590 2732.810 219.770 ;
        RECT 2733.230 218.590 2734.410 219.770 ;
        RECT 2731.630 216.990 2732.810 218.170 ;
        RECT 2733.230 216.990 2734.410 218.170 ;
        RECT 2731.630 38.590 2732.810 39.770 ;
        RECT 2733.230 38.590 2734.410 39.770 ;
        RECT 2731.630 36.990 2732.810 38.170 ;
        RECT 2733.230 36.990 2734.410 38.170 ;
        RECT 2731.630 -9.260 2732.810 -8.080 ;
        RECT 2733.230 -9.260 2734.410 -8.080 ;
        RECT 2731.630 -10.860 2732.810 -9.680 ;
        RECT 2733.230 -10.860 2734.410 -9.680 ;
        RECT 2911.630 3529.360 2912.810 3530.540 ;
        RECT 2913.230 3529.360 2914.410 3530.540 ;
        RECT 2911.630 3527.760 2912.810 3528.940 ;
        RECT 2913.230 3527.760 2914.410 3528.940 ;
        RECT 2911.630 3458.590 2912.810 3459.770 ;
        RECT 2913.230 3458.590 2914.410 3459.770 ;
        RECT 2911.630 3456.990 2912.810 3458.170 ;
        RECT 2913.230 3456.990 2914.410 3458.170 ;
        RECT 2911.630 3278.590 2912.810 3279.770 ;
        RECT 2913.230 3278.590 2914.410 3279.770 ;
        RECT 2911.630 3276.990 2912.810 3278.170 ;
        RECT 2913.230 3276.990 2914.410 3278.170 ;
        RECT 2911.630 3098.590 2912.810 3099.770 ;
        RECT 2913.230 3098.590 2914.410 3099.770 ;
        RECT 2911.630 3096.990 2912.810 3098.170 ;
        RECT 2913.230 3096.990 2914.410 3098.170 ;
        RECT 2911.630 2918.590 2912.810 2919.770 ;
        RECT 2913.230 2918.590 2914.410 2919.770 ;
        RECT 2911.630 2916.990 2912.810 2918.170 ;
        RECT 2913.230 2916.990 2914.410 2918.170 ;
        RECT 2911.630 2738.590 2912.810 2739.770 ;
        RECT 2913.230 2738.590 2914.410 2739.770 ;
        RECT 2911.630 2736.990 2912.810 2738.170 ;
        RECT 2913.230 2736.990 2914.410 2738.170 ;
        RECT 2911.630 2558.590 2912.810 2559.770 ;
        RECT 2913.230 2558.590 2914.410 2559.770 ;
        RECT 2911.630 2556.990 2912.810 2558.170 ;
        RECT 2913.230 2556.990 2914.410 2558.170 ;
        RECT 2911.630 2378.590 2912.810 2379.770 ;
        RECT 2913.230 2378.590 2914.410 2379.770 ;
        RECT 2911.630 2376.990 2912.810 2378.170 ;
        RECT 2913.230 2376.990 2914.410 2378.170 ;
        RECT 2911.630 2198.590 2912.810 2199.770 ;
        RECT 2913.230 2198.590 2914.410 2199.770 ;
        RECT 2911.630 2196.990 2912.810 2198.170 ;
        RECT 2913.230 2196.990 2914.410 2198.170 ;
        RECT 2911.630 2018.590 2912.810 2019.770 ;
        RECT 2913.230 2018.590 2914.410 2019.770 ;
        RECT 2911.630 2016.990 2912.810 2018.170 ;
        RECT 2913.230 2016.990 2914.410 2018.170 ;
        RECT 2911.630 1838.590 2912.810 1839.770 ;
        RECT 2913.230 1838.590 2914.410 1839.770 ;
        RECT 2911.630 1836.990 2912.810 1838.170 ;
        RECT 2913.230 1836.990 2914.410 1838.170 ;
        RECT 2911.630 1658.590 2912.810 1659.770 ;
        RECT 2913.230 1658.590 2914.410 1659.770 ;
        RECT 2911.630 1656.990 2912.810 1658.170 ;
        RECT 2913.230 1656.990 2914.410 1658.170 ;
        RECT 2911.630 1478.590 2912.810 1479.770 ;
        RECT 2913.230 1478.590 2914.410 1479.770 ;
        RECT 2911.630 1476.990 2912.810 1478.170 ;
        RECT 2913.230 1476.990 2914.410 1478.170 ;
        RECT 2911.630 1298.590 2912.810 1299.770 ;
        RECT 2913.230 1298.590 2914.410 1299.770 ;
        RECT 2911.630 1296.990 2912.810 1298.170 ;
        RECT 2913.230 1296.990 2914.410 1298.170 ;
        RECT 2911.630 1118.590 2912.810 1119.770 ;
        RECT 2913.230 1118.590 2914.410 1119.770 ;
        RECT 2911.630 1116.990 2912.810 1118.170 ;
        RECT 2913.230 1116.990 2914.410 1118.170 ;
        RECT 2911.630 938.590 2912.810 939.770 ;
        RECT 2913.230 938.590 2914.410 939.770 ;
        RECT 2911.630 936.990 2912.810 938.170 ;
        RECT 2913.230 936.990 2914.410 938.170 ;
        RECT 2911.630 758.590 2912.810 759.770 ;
        RECT 2913.230 758.590 2914.410 759.770 ;
        RECT 2911.630 756.990 2912.810 758.170 ;
        RECT 2913.230 756.990 2914.410 758.170 ;
        RECT 2911.630 578.590 2912.810 579.770 ;
        RECT 2913.230 578.590 2914.410 579.770 ;
        RECT 2911.630 576.990 2912.810 578.170 ;
        RECT 2913.230 576.990 2914.410 578.170 ;
        RECT 2911.630 398.590 2912.810 399.770 ;
        RECT 2913.230 398.590 2914.410 399.770 ;
        RECT 2911.630 396.990 2912.810 398.170 ;
        RECT 2913.230 396.990 2914.410 398.170 ;
        RECT 2911.630 218.590 2912.810 219.770 ;
        RECT 2913.230 218.590 2914.410 219.770 ;
        RECT 2911.630 216.990 2912.810 218.170 ;
        RECT 2913.230 216.990 2914.410 218.170 ;
        RECT 2911.630 38.590 2912.810 39.770 ;
        RECT 2913.230 38.590 2914.410 39.770 ;
        RECT 2911.630 36.990 2912.810 38.170 ;
        RECT 2913.230 36.990 2914.410 38.170 ;
        RECT 2911.630 -9.260 2912.810 -8.080 ;
        RECT 2913.230 -9.260 2914.410 -8.080 ;
        RECT 2911.630 -10.860 2912.810 -9.680 ;
        RECT 2913.230 -10.860 2914.410 -9.680 ;
        RECT 2933.060 3529.360 2934.240 3530.540 ;
        RECT 2934.660 3529.360 2935.840 3530.540 ;
        RECT 2933.060 3527.760 2934.240 3528.940 ;
        RECT 2934.660 3527.760 2935.840 3528.940 ;
        RECT 2933.060 3458.590 2934.240 3459.770 ;
        RECT 2934.660 3458.590 2935.840 3459.770 ;
        RECT 2933.060 3456.990 2934.240 3458.170 ;
        RECT 2934.660 3456.990 2935.840 3458.170 ;
        RECT 2933.060 3278.590 2934.240 3279.770 ;
        RECT 2934.660 3278.590 2935.840 3279.770 ;
        RECT 2933.060 3276.990 2934.240 3278.170 ;
        RECT 2934.660 3276.990 2935.840 3278.170 ;
        RECT 2933.060 3098.590 2934.240 3099.770 ;
        RECT 2934.660 3098.590 2935.840 3099.770 ;
        RECT 2933.060 3096.990 2934.240 3098.170 ;
        RECT 2934.660 3096.990 2935.840 3098.170 ;
        RECT 2933.060 2918.590 2934.240 2919.770 ;
        RECT 2934.660 2918.590 2935.840 2919.770 ;
        RECT 2933.060 2916.990 2934.240 2918.170 ;
        RECT 2934.660 2916.990 2935.840 2918.170 ;
        RECT 2933.060 2738.590 2934.240 2739.770 ;
        RECT 2934.660 2738.590 2935.840 2739.770 ;
        RECT 2933.060 2736.990 2934.240 2738.170 ;
        RECT 2934.660 2736.990 2935.840 2738.170 ;
        RECT 2933.060 2558.590 2934.240 2559.770 ;
        RECT 2934.660 2558.590 2935.840 2559.770 ;
        RECT 2933.060 2556.990 2934.240 2558.170 ;
        RECT 2934.660 2556.990 2935.840 2558.170 ;
        RECT 2933.060 2378.590 2934.240 2379.770 ;
        RECT 2934.660 2378.590 2935.840 2379.770 ;
        RECT 2933.060 2376.990 2934.240 2378.170 ;
        RECT 2934.660 2376.990 2935.840 2378.170 ;
        RECT 2933.060 2198.590 2934.240 2199.770 ;
        RECT 2934.660 2198.590 2935.840 2199.770 ;
        RECT 2933.060 2196.990 2934.240 2198.170 ;
        RECT 2934.660 2196.990 2935.840 2198.170 ;
        RECT 2933.060 2018.590 2934.240 2019.770 ;
        RECT 2934.660 2018.590 2935.840 2019.770 ;
        RECT 2933.060 2016.990 2934.240 2018.170 ;
        RECT 2934.660 2016.990 2935.840 2018.170 ;
        RECT 2933.060 1838.590 2934.240 1839.770 ;
        RECT 2934.660 1838.590 2935.840 1839.770 ;
        RECT 2933.060 1836.990 2934.240 1838.170 ;
        RECT 2934.660 1836.990 2935.840 1838.170 ;
        RECT 2933.060 1658.590 2934.240 1659.770 ;
        RECT 2934.660 1658.590 2935.840 1659.770 ;
        RECT 2933.060 1656.990 2934.240 1658.170 ;
        RECT 2934.660 1656.990 2935.840 1658.170 ;
        RECT 2933.060 1478.590 2934.240 1479.770 ;
        RECT 2934.660 1478.590 2935.840 1479.770 ;
        RECT 2933.060 1476.990 2934.240 1478.170 ;
        RECT 2934.660 1476.990 2935.840 1478.170 ;
        RECT 2933.060 1298.590 2934.240 1299.770 ;
        RECT 2934.660 1298.590 2935.840 1299.770 ;
        RECT 2933.060 1296.990 2934.240 1298.170 ;
        RECT 2934.660 1296.990 2935.840 1298.170 ;
        RECT 2933.060 1118.590 2934.240 1119.770 ;
        RECT 2934.660 1118.590 2935.840 1119.770 ;
        RECT 2933.060 1116.990 2934.240 1118.170 ;
        RECT 2934.660 1116.990 2935.840 1118.170 ;
        RECT 2933.060 938.590 2934.240 939.770 ;
        RECT 2934.660 938.590 2935.840 939.770 ;
        RECT 2933.060 936.990 2934.240 938.170 ;
        RECT 2934.660 936.990 2935.840 938.170 ;
        RECT 2933.060 758.590 2934.240 759.770 ;
        RECT 2934.660 758.590 2935.840 759.770 ;
        RECT 2933.060 756.990 2934.240 758.170 ;
        RECT 2934.660 756.990 2935.840 758.170 ;
        RECT 2933.060 578.590 2934.240 579.770 ;
        RECT 2934.660 578.590 2935.840 579.770 ;
        RECT 2933.060 576.990 2934.240 578.170 ;
        RECT 2934.660 576.990 2935.840 578.170 ;
        RECT 2933.060 398.590 2934.240 399.770 ;
        RECT 2934.660 398.590 2935.840 399.770 ;
        RECT 2933.060 396.990 2934.240 398.170 ;
        RECT 2934.660 396.990 2935.840 398.170 ;
        RECT 2933.060 218.590 2934.240 219.770 ;
        RECT 2934.660 218.590 2935.840 219.770 ;
        RECT 2933.060 216.990 2934.240 218.170 ;
        RECT 2934.660 216.990 2935.840 218.170 ;
        RECT 2933.060 38.590 2934.240 39.770 ;
        RECT 2934.660 38.590 2935.840 39.770 ;
        RECT 2933.060 36.990 2934.240 38.170 ;
        RECT 2934.660 36.990 2935.840 38.170 ;
        RECT 2933.060 -9.260 2934.240 -8.080 ;
        RECT 2934.660 -9.260 2935.840 -8.080 ;
        RECT 2933.060 -10.860 2934.240 -9.680 ;
        RECT 2934.660 -10.860 2935.840 -9.680 ;
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
        RECT -45.180 3456.830 2964.800 3459.930 ;
        RECT -45.180 3276.830 2964.800 3279.930 ;
        RECT -45.180 3096.830 2964.800 3099.930 ;
        RECT -45.180 2916.830 2964.800 2919.930 ;
        RECT -45.180 2736.830 2964.800 2739.930 ;
        RECT -45.180 2556.830 2964.800 2559.930 ;
        RECT -45.180 2376.830 2964.800 2379.930 ;
        RECT -45.180 2196.830 2964.800 2199.930 ;
        RECT -45.180 2016.830 2964.800 2019.930 ;
        RECT -45.180 1836.830 2964.800 1839.930 ;
        RECT -45.180 1656.830 2964.800 1659.930 ;
        RECT -45.180 1476.830 2964.800 1479.930 ;
        RECT -45.180 1296.830 2964.800 1299.930 ;
        RECT -45.180 1116.830 2964.800 1119.930 ;
        RECT -45.180 936.830 2964.800 939.930 ;
        RECT -45.180 756.830 2964.800 759.930 ;
        RECT -45.180 576.830 2964.800 579.930 ;
        RECT -45.180 396.830 2964.800 399.930 ;
        RECT -45.180 216.830 2964.800 219.930 ;
        RECT -45.180 36.830 2964.800 39.930 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -25.980 -20.620 -22.880 3540.300 ;
        RECT 76.470 -39.820 79.570 3559.500 ;
        RECT 256.470 -39.820 259.570 3559.500 ;
        RECT 436.470 760.000 439.570 3559.500 ;
        RECT 616.470 760.000 619.570 3559.500 ;
        RECT 436.470 -39.820 439.570 490.000 ;
        RECT 616.470 -39.820 619.570 490.000 ;
        RECT 796.470 -39.820 799.570 3559.500 ;
        RECT 976.470 -39.820 979.570 3559.500 ;
        RECT 1156.470 -39.820 1159.570 3559.500 ;
        RECT 1336.470 -39.820 1339.570 3559.500 ;
        RECT 1516.470 -39.820 1519.570 3559.500 ;
        RECT 1696.470 -39.820 1699.570 3559.500 ;
        RECT 1876.470 -39.820 1879.570 3559.500 ;
        RECT 2056.470 -39.820 2059.570 3559.500 ;
        RECT 2236.470 -39.820 2239.570 3559.500 ;
        RECT 2416.470 -39.820 2419.570 3559.500 ;
        RECT 2596.470 -39.820 2599.570 3559.500 ;
        RECT 2776.470 -39.820 2779.570 3559.500 ;
        RECT 2942.500 -20.620 2945.600 3540.300 ;
      LAYER via4 ;
        RECT -25.820 3538.960 -24.640 3540.140 ;
        RECT -24.220 3538.960 -23.040 3540.140 ;
        RECT -25.820 3537.360 -24.640 3538.540 ;
        RECT -24.220 3537.360 -23.040 3538.540 ;
        RECT -25.820 3503.590 -24.640 3504.770 ;
        RECT -24.220 3503.590 -23.040 3504.770 ;
        RECT -25.820 3501.990 -24.640 3503.170 ;
        RECT -24.220 3501.990 -23.040 3503.170 ;
        RECT -25.820 3323.590 -24.640 3324.770 ;
        RECT -24.220 3323.590 -23.040 3324.770 ;
        RECT -25.820 3321.990 -24.640 3323.170 ;
        RECT -24.220 3321.990 -23.040 3323.170 ;
        RECT -25.820 3143.590 -24.640 3144.770 ;
        RECT -24.220 3143.590 -23.040 3144.770 ;
        RECT -25.820 3141.990 -24.640 3143.170 ;
        RECT -24.220 3141.990 -23.040 3143.170 ;
        RECT -25.820 2963.590 -24.640 2964.770 ;
        RECT -24.220 2963.590 -23.040 2964.770 ;
        RECT -25.820 2961.990 -24.640 2963.170 ;
        RECT -24.220 2961.990 -23.040 2963.170 ;
        RECT -25.820 2783.590 -24.640 2784.770 ;
        RECT -24.220 2783.590 -23.040 2784.770 ;
        RECT -25.820 2781.990 -24.640 2783.170 ;
        RECT -24.220 2781.990 -23.040 2783.170 ;
        RECT -25.820 2603.590 -24.640 2604.770 ;
        RECT -24.220 2603.590 -23.040 2604.770 ;
        RECT -25.820 2601.990 -24.640 2603.170 ;
        RECT -24.220 2601.990 -23.040 2603.170 ;
        RECT -25.820 2423.590 -24.640 2424.770 ;
        RECT -24.220 2423.590 -23.040 2424.770 ;
        RECT -25.820 2421.990 -24.640 2423.170 ;
        RECT -24.220 2421.990 -23.040 2423.170 ;
        RECT -25.820 2243.590 -24.640 2244.770 ;
        RECT -24.220 2243.590 -23.040 2244.770 ;
        RECT -25.820 2241.990 -24.640 2243.170 ;
        RECT -24.220 2241.990 -23.040 2243.170 ;
        RECT -25.820 2063.590 -24.640 2064.770 ;
        RECT -24.220 2063.590 -23.040 2064.770 ;
        RECT -25.820 2061.990 -24.640 2063.170 ;
        RECT -24.220 2061.990 -23.040 2063.170 ;
        RECT -25.820 1883.590 -24.640 1884.770 ;
        RECT -24.220 1883.590 -23.040 1884.770 ;
        RECT -25.820 1881.990 -24.640 1883.170 ;
        RECT -24.220 1881.990 -23.040 1883.170 ;
        RECT -25.820 1703.590 -24.640 1704.770 ;
        RECT -24.220 1703.590 -23.040 1704.770 ;
        RECT -25.820 1701.990 -24.640 1703.170 ;
        RECT -24.220 1701.990 -23.040 1703.170 ;
        RECT -25.820 1523.590 -24.640 1524.770 ;
        RECT -24.220 1523.590 -23.040 1524.770 ;
        RECT -25.820 1521.990 -24.640 1523.170 ;
        RECT -24.220 1521.990 -23.040 1523.170 ;
        RECT -25.820 1343.590 -24.640 1344.770 ;
        RECT -24.220 1343.590 -23.040 1344.770 ;
        RECT -25.820 1341.990 -24.640 1343.170 ;
        RECT -24.220 1341.990 -23.040 1343.170 ;
        RECT -25.820 1163.590 -24.640 1164.770 ;
        RECT -24.220 1163.590 -23.040 1164.770 ;
        RECT -25.820 1161.990 -24.640 1163.170 ;
        RECT -24.220 1161.990 -23.040 1163.170 ;
        RECT -25.820 983.590 -24.640 984.770 ;
        RECT -24.220 983.590 -23.040 984.770 ;
        RECT -25.820 981.990 -24.640 983.170 ;
        RECT -24.220 981.990 -23.040 983.170 ;
        RECT -25.820 803.590 -24.640 804.770 ;
        RECT -24.220 803.590 -23.040 804.770 ;
        RECT -25.820 801.990 -24.640 803.170 ;
        RECT -24.220 801.990 -23.040 803.170 ;
        RECT -25.820 623.590 -24.640 624.770 ;
        RECT -24.220 623.590 -23.040 624.770 ;
        RECT -25.820 621.990 -24.640 623.170 ;
        RECT -24.220 621.990 -23.040 623.170 ;
        RECT -25.820 443.590 -24.640 444.770 ;
        RECT -24.220 443.590 -23.040 444.770 ;
        RECT -25.820 441.990 -24.640 443.170 ;
        RECT -24.220 441.990 -23.040 443.170 ;
        RECT -25.820 263.590 -24.640 264.770 ;
        RECT -24.220 263.590 -23.040 264.770 ;
        RECT -25.820 261.990 -24.640 263.170 ;
        RECT -24.220 261.990 -23.040 263.170 ;
        RECT -25.820 83.590 -24.640 84.770 ;
        RECT -24.220 83.590 -23.040 84.770 ;
        RECT -25.820 81.990 -24.640 83.170 ;
        RECT -24.220 81.990 -23.040 83.170 ;
        RECT -25.820 -18.860 -24.640 -17.680 ;
        RECT -24.220 -18.860 -23.040 -17.680 ;
        RECT -25.820 -20.460 -24.640 -19.280 ;
        RECT -24.220 -20.460 -23.040 -19.280 ;
        RECT 76.630 3538.960 77.810 3540.140 ;
        RECT 78.230 3538.960 79.410 3540.140 ;
        RECT 76.630 3537.360 77.810 3538.540 ;
        RECT 78.230 3537.360 79.410 3538.540 ;
        RECT 76.630 3503.590 77.810 3504.770 ;
        RECT 78.230 3503.590 79.410 3504.770 ;
        RECT 76.630 3501.990 77.810 3503.170 ;
        RECT 78.230 3501.990 79.410 3503.170 ;
        RECT 76.630 3323.590 77.810 3324.770 ;
        RECT 78.230 3323.590 79.410 3324.770 ;
        RECT 76.630 3321.990 77.810 3323.170 ;
        RECT 78.230 3321.990 79.410 3323.170 ;
        RECT 76.630 3143.590 77.810 3144.770 ;
        RECT 78.230 3143.590 79.410 3144.770 ;
        RECT 76.630 3141.990 77.810 3143.170 ;
        RECT 78.230 3141.990 79.410 3143.170 ;
        RECT 76.630 2963.590 77.810 2964.770 ;
        RECT 78.230 2963.590 79.410 2964.770 ;
        RECT 76.630 2961.990 77.810 2963.170 ;
        RECT 78.230 2961.990 79.410 2963.170 ;
        RECT 76.630 2783.590 77.810 2784.770 ;
        RECT 78.230 2783.590 79.410 2784.770 ;
        RECT 76.630 2781.990 77.810 2783.170 ;
        RECT 78.230 2781.990 79.410 2783.170 ;
        RECT 76.630 2603.590 77.810 2604.770 ;
        RECT 78.230 2603.590 79.410 2604.770 ;
        RECT 76.630 2601.990 77.810 2603.170 ;
        RECT 78.230 2601.990 79.410 2603.170 ;
        RECT 76.630 2423.590 77.810 2424.770 ;
        RECT 78.230 2423.590 79.410 2424.770 ;
        RECT 76.630 2421.990 77.810 2423.170 ;
        RECT 78.230 2421.990 79.410 2423.170 ;
        RECT 76.630 2243.590 77.810 2244.770 ;
        RECT 78.230 2243.590 79.410 2244.770 ;
        RECT 76.630 2241.990 77.810 2243.170 ;
        RECT 78.230 2241.990 79.410 2243.170 ;
        RECT 76.630 2063.590 77.810 2064.770 ;
        RECT 78.230 2063.590 79.410 2064.770 ;
        RECT 76.630 2061.990 77.810 2063.170 ;
        RECT 78.230 2061.990 79.410 2063.170 ;
        RECT 76.630 1883.590 77.810 1884.770 ;
        RECT 78.230 1883.590 79.410 1884.770 ;
        RECT 76.630 1881.990 77.810 1883.170 ;
        RECT 78.230 1881.990 79.410 1883.170 ;
        RECT 76.630 1703.590 77.810 1704.770 ;
        RECT 78.230 1703.590 79.410 1704.770 ;
        RECT 76.630 1701.990 77.810 1703.170 ;
        RECT 78.230 1701.990 79.410 1703.170 ;
        RECT 76.630 1523.590 77.810 1524.770 ;
        RECT 78.230 1523.590 79.410 1524.770 ;
        RECT 76.630 1521.990 77.810 1523.170 ;
        RECT 78.230 1521.990 79.410 1523.170 ;
        RECT 76.630 1343.590 77.810 1344.770 ;
        RECT 78.230 1343.590 79.410 1344.770 ;
        RECT 76.630 1341.990 77.810 1343.170 ;
        RECT 78.230 1341.990 79.410 1343.170 ;
        RECT 76.630 1163.590 77.810 1164.770 ;
        RECT 78.230 1163.590 79.410 1164.770 ;
        RECT 76.630 1161.990 77.810 1163.170 ;
        RECT 78.230 1161.990 79.410 1163.170 ;
        RECT 76.630 983.590 77.810 984.770 ;
        RECT 78.230 983.590 79.410 984.770 ;
        RECT 76.630 981.990 77.810 983.170 ;
        RECT 78.230 981.990 79.410 983.170 ;
        RECT 76.630 803.590 77.810 804.770 ;
        RECT 78.230 803.590 79.410 804.770 ;
        RECT 76.630 801.990 77.810 803.170 ;
        RECT 78.230 801.990 79.410 803.170 ;
        RECT 76.630 623.590 77.810 624.770 ;
        RECT 78.230 623.590 79.410 624.770 ;
        RECT 76.630 621.990 77.810 623.170 ;
        RECT 78.230 621.990 79.410 623.170 ;
        RECT 76.630 443.590 77.810 444.770 ;
        RECT 78.230 443.590 79.410 444.770 ;
        RECT 76.630 441.990 77.810 443.170 ;
        RECT 78.230 441.990 79.410 443.170 ;
        RECT 76.630 263.590 77.810 264.770 ;
        RECT 78.230 263.590 79.410 264.770 ;
        RECT 76.630 261.990 77.810 263.170 ;
        RECT 78.230 261.990 79.410 263.170 ;
        RECT 76.630 83.590 77.810 84.770 ;
        RECT 78.230 83.590 79.410 84.770 ;
        RECT 76.630 81.990 77.810 83.170 ;
        RECT 78.230 81.990 79.410 83.170 ;
        RECT 76.630 -18.860 77.810 -17.680 ;
        RECT 78.230 -18.860 79.410 -17.680 ;
        RECT 76.630 -20.460 77.810 -19.280 ;
        RECT 78.230 -20.460 79.410 -19.280 ;
        RECT 256.630 3538.960 257.810 3540.140 ;
        RECT 258.230 3538.960 259.410 3540.140 ;
        RECT 256.630 3537.360 257.810 3538.540 ;
        RECT 258.230 3537.360 259.410 3538.540 ;
        RECT 256.630 3503.590 257.810 3504.770 ;
        RECT 258.230 3503.590 259.410 3504.770 ;
        RECT 256.630 3501.990 257.810 3503.170 ;
        RECT 258.230 3501.990 259.410 3503.170 ;
        RECT 256.630 3323.590 257.810 3324.770 ;
        RECT 258.230 3323.590 259.410 3324.770 ;
        RECT 256.630 3321.990 257.810 3323.170 ;
        RECT 258.230 3321.990 259.410 3323.170 ;
        RECT 256.630 3143.590 257.810 3144.770 ;
        RECT 258.230 3143.590 259.410 3144.770 ;
        RECT 256.630 3141.990 257.810 3143.170 ;
        RECT 258.230 3141.990 259.410 3143.170 ;
        RECT 256.630 2963.590 257.810 2964.770 ;
        RECT 258.230 2963.590 259.410 2964.770 ;
        RECT 256.630 2961.990 257.810 2963.170 ;
        RECT 258.230 2961.990 259.410 2963.170 ;
        RECT 256.630 2783.590 257.810 2784.770 ;
        RECT 258.230 2783.590 259.410 2784.770 ;
        RECT 256.630 2781.990 257.810 2783.170 ;
        RECT 258.230 2781.990 259.410 2783.170 ;
        RECT 256.630 2603.590 257.810 2604.770 ;
        RECT 258.230 2603.590 259.410 2604.770 ;
        RECT 256.630 2601.990 257.810 2603.170 ;
        RECT 258.230 2601.990 259.410 2603.170 ;
        RECT 256.630 2423.590 257.810 2424.770 ;
        RECT 258.230 2423.590 259.410 2424.770 ;
        RECT 256.630 2421.990 257.810 2423.170 ;
        RECT 258.230 2421.990 259.410 2423.170 ;
        RECT 256.630 2243.590 257.810 2244.770 ;
        RECT 258.230 2243.590 259.410 2244.770 ;
        RECT 256.630 2241.990 257.810 2243.170 ;
        RECT 258.230 2241.990 259.410 2243.170 ;
        RECT 256.630 2063.590 257.810 2064.770 ;
        RECT 258.230 2063.590 259.410 2064.770 ;
        RECT 256.630 2061.990 257.810 2063.170 ;
        RECT 258.230 2061.990 259.410 2063.170 ;
        RECT 256.630 1883.590 257.810 1884.770 ;
        RECT 258.230 1883.590 259.410 1884.770 ;
        RECT 256.630 1881.990 257.810 1883.170 ;
        RECT 258.230 1881.990 259.410 1883.170 ;
        RECT 256.630 1703.590 257.810 1704.770 ;
        RECT 258.230 1703.590 259.410 1704.770 ;
        RECT 256.630 1701.990 257.810 1703.170 ;
        RECT 258.230 1701.990 259.410 1703.170 ;
        RECT 256.630 1523.590 257.810 1524.770 ;
        RECT 258.230 1523.590 259.410 1524.770 ;
        RECT 256.630 1521.990 257.810 1523.170 ;
        RECT 258.230 1521.990 259.410 1523.170 ;
        RECT 256.630 1343.590 257.810 1344.770 ;
        RECT 258.230 1343.590 259.410 1344.770 ;
        RECT 256.630 1341.990 257.810 1343.170 ;
        RECT 258.230 1341.990 259.410 1343.170 ;
        RECT 256.630 1163.590 257.810 1164.770 ;
        RECT 258.230 1163.590 259.410 1164.770 ;
        RECT 256.630 1161.990 257.810 1163.170 ;
        RECT 258.230 1161.990 259.410 1163.170 ;
        RECT 256.630 983.590 257.810 984.770 ;
        RECT 258.230 983.590 259.410 984.770 ;
        RECT 256.630 981.990 257.810 983.170 ;
        RECT 258.230 981.990 259.410 983.170 ;
        RECT 256.630 803.590 257.810 804.770 ;
        RECT 258.230 803.590 259.410 804.770 ;
        RECT 256.630 801.990 257.810 803.170 ;
        RECT 258.230 801.990 259.410 803.170 ;
        RECT 436.630 3538.960 437.810 3540.140 ;
        RECT 438.230 3538.960 439.410 3540.140 ;
        RECT 436.630 3537.360 437.810 3538.540 ;
        RECT 438.230 3537.360 439.410 3538.540 ;
        RECT 436.630 3503.590 437.810 3504.770 ;
        RECT 438.230 3503.590 439.410 3504.770 ;
        RECT 436.630 3501.990 437.810 3503.170 ;
        RECT 438.230 3501.990 439.410 3503.170 ;
        RECT 436.630 3323.590 437.810 3324.770 ;
        RECT 438.230 3323.590 439.410 3324.770 ;
        RECT 436.630 3321.990 437.810 3323.170 ;
        RECT 438.230 3321.990 439.410 3323.170 ;
        RECT 436.630 3143.590 437.810 3144.770 ;
        RECT 438.230 3143.590 439.410 3144.770 ;
        RECT 436.630 3141.990 437.810 3143.170 ;
        RECT 438.230 3141.990 439.410 3143.170 ;
        RECT 436.630 2963.590 437.810 2964.770 ;
        RECT 438.230 2963.590 439.410 2964.770 ;
        RECT 436.630 2961.990 437.810 2963.170 ;
        RECT 438.230 2961.990 439.410 2963.170 ;
        RECT 436.630 2783.590 437.810 2784.770 ;
        RECT 438.230 2783.590 439.410 2784.770 ;
        RECT 436.630 2781.990 437.810 2783.170 ;
        RECT 438.230 2781.990 439.410 2783.170 ;
        RECT 436.630 2603.590 437.810 2604.770 ;
        RECT 438.230 2603.590 439.410 2604.770 ;
        RECT 436.630 2601.990 437.810 2603.170 ;
        RECT 438.230 2601.990 439.410 2603.170 ;
        RECT 436.630 2423.590 437.810 2424.770 ;
        RECT 438.230 2423.590 439.410 2424.770 ;
        RECT 436.630 2421.990 437.810 2423.170 ;
        RECT 438.230 2421.990 439.410 2423.170 ;
        RECT 436.630 2243.590 437.810 2244.770 ;
        RECT 438.230 2243.590 439.410 2244.770 ;
        RECT 436.630 2241.990 437.810 2243.170 ;
        RECT 438.230 2241.990 439.410 2243.170 ;
        RECT 436.630 2063.590 437.810 2064.770 ;
        RECT 438.230 2063.590 439.410 2064.770 ;
        RECT 436.630 2061.990 437.810 2063.170 ;
        RECT 438.230 2061.990 439.410 2063.170 ;
        RECT 436.630 1883.590 437.810 1884.770 ;
        RECT 438.230 1883.590 439.410 1884.770 ;
        RECT 436.630 1881.990 437.810 1883.170 ;
        RECT 438.230 1881.990 439.410 1883.170 ;
        RECT 436.630 1703.590 437.810 1704.770 ;
        RECT 438.230 1703.590 439.410 1704.770 ;
        RECT 436.630 1701.990 437.810 1703.170 ;
        RECT 438.230 1701.990 439.410 1703.170 ;
        RECT 436.630 1523.590 437.810 1524.770 ;
        RECT 438.230 1523.590 439.410 1524.770 ;
        RECT 436.630 1521.990 437.810 1523.170 ;
        RECT 438.230 1521.990 439.410 1523.170 ;
        RECT 436.630 1343.590 437.810 1344.770 ;
        RECT 438.230 1343.590 439.410 1344.770 ;
        RECT 436.630 1341.990 437.810 1343.170 ;
        RECT 438.230 1341.990 439.410 1343.170 ;
        RECT 436.630 1163.590 437.810 1164.770 ;
        RECT 438.230 1163.590 439.410 1164.770 ;
        RECT 436.630 1161.990 437.810 1163.170 ;
        RECT 438.230 1161.990 439.410 1163.170 ;
        RECT 436.630 983.590 437.810 984.770 ;
        RECT 438.230 983.590 439.410 984.770 ;
        RECT 436.630 981.990 437.810 983.170 ;
        RECT 438.230 981.990 439.410 983.170 ;
        RECT 436.630 803.590 437.810 804.770 ;
        RECT 438.230 803.590 439.410 804.770 ;
        RECT 436.630 801.990 437.810 803.170 ;
        RECT 438.230 801.990 439.410 803.170 ;
        RECT 616.630 3538.960 617.810 3540.140 ;
        RECT 618.230 3538.960 619.410 3540.140 ;
        RECT 616.630 3537.360 617.810 3538.540 ;
        RECT 618.230 3537.360 619.410 3538.540 ;
        RECT 616.630 3503.590 617.810 3504.770 ;
        RECT 618.230 3503.590 619.410 3504.770 ;
        RECT 616.630 3501.990 617.810 3503.170 ;
        RECT 618.230 3501.990 619.410 3503.170 ;
        RECT 616.630 3323.590 617.810 3324.770 ;
        RECT 618.230 3323.590 619.410 3324.770 ;
        RECT 616.630 3321.990 617.810 3323.170 ;
        RECT 618.230 3321.990 619.410 3323.170 ;
        RECT 616.630 3143.590 617.810 3144.770 ;
        RECT 618.230 3143.590 619.410 3144.770 ;
        RECT 616.630 3141.990 617.810 3143.170 ;
        RECT 618.230 3141.990 619.410 3143.170 ;
        RECT 616.630 2963.590 617.810 2964.770 ;
        RECT 618.230 2963.590 619.410 2964.770 ;
        RECT 616.630 2961.990 617.810 2963.170 ;
        RECT 618.230 2961.990 619.410 2963.170 ;
        RECT 616.630 2783.590 617.810 2784.770 ;
        RECT 618.230 2783.590 619.410 2784.770 ;
        RECT 616.630 2781.990 617.810 2783.170 ;
        RECT 618.230 2781.990 619.410 2783.170 ;
        RECT 616.630 2603.590 617.810 2604.770 ;
        RECT 618.230 2603.590 619.410 2604.770 ;
        RECT 616.630 2601.990 617.810 2603.170 ;
        RECT 618.230 2601.990 619.410 2603.170 ;
        RECT 616.630 2423.590 617.810 2424.770 ;
        RECT 618.230 2423.590 619.410 2424.770 ;
        RECT 616.630 2421.990 617.810 2423.170 ;
        RECT 618.230 2421.990 619.410 2423.170 ;
        RECT 616.630 2243.590 617.810 2244.770 ;
        RECT 618.230 2243.590 619.410 2244.770 ;
        RECT 616.630 2241.990 617.810 2243.170 ;
        RECT 618.230 2241.990 619.410 2243.170 ;
        RECT 616.630 2063.590 617.810 2064.770 ;
        RECT 618.230 2063.590 619.410 2064.770 ;
        RECT 616.630 2061.990 617.810 2063.170 ;
        RECT 618.230 2061.990 619.410 2063.170 ;
        RECT 616.630 1883.590 617.810 1884.770 ;
        RECT 618.230 1883.590 619.410 1884.770 ;
        RECT 616.630 1881.990 617.810 1883.170 ;
        RECT 618.230 1881.990 619.410 1883.170 ;
        RECT 616.630 1703.590 617.810 1704.770 ;
        RECT 618.230 1703.590 619.410 1704.770 ;
        RECT 616.630 1701.990 617.810 1703.170 ;
        RECT 618.230 1701.990 619.410 1703.170 ;
        RECT 616.630 1523.590 617.810 1524.770 ;
        RECT 618.230 1523.590 619.410 1524.770 ;
        RECT 616.630 1521.990 617.810 1523.170 ;
        RECT 618.230 1521.990 619.410 1523.170 ;
        RECT 616.630 1343.590 617.810 1344.770 ;
        RECT 618.230 1343.590 619.410 1344.770 ;
        RECT 616.630 1341.990 617.810 1343.170 ;
        RECT 618.230 1341.990 619.410 1343.170 ;
        RECT 616.630 1163.590 617.810 1164.770 ;
        RECT 618.230 1163.590 619.410 1164.770 ;
        RECT 616.630 1161.990 617.810 1163.170 ;
        RECT 618.230 1161.990 619.410 1163.170 ;
        RECT 616.630 983.590 617.810 984.770 ;
        RECT 618.230 983.590 619.410 984.770 ;
        RECT 616.630 981.990 617.810 983.170 ;
        RECT 618.230 981.990 619.410 983.170 ;
        RECT 616.630 803.590 617.810 804.770 ;
        RECT 618.230 803.590 619.410 804.770 ;
        RECT 616.630 801.990 617.810 803.170 ;
        RECT 618.230 801.990 619.410 803.170 ;
        RECT 796.630 3538.960 797.810 3540.140 ;
        RECT 798.230 3538.960 799.410 3540.140 ;
        RECT 796.630 3537.360 797.810 3538.540 ;
        RECT 798.230 3537.360 799.410 3538.540 ;
        RECT 796.630 3503.590 797.810 3504.770 ;
        RECT 798.230 3503.590 799.410 3504.770 ;
        RECT 796.630 3501.990 797.810 3503.170 ;
        RECT 798.230 3501.990 799.410 3503.170 ;
        RECT 796.630 3323.590 797.810 3324.770 ;
        RECT 798.230 3323.590 799.410 3324.770 ;
        RECT 796.630 3321.990 797.810 3323.170 ;
        RECT 798.230 3321.990 799.410 3323.170 ;
        RECT 796.630 3143.590 797.810 3144.770 ;
        RECT 798.230 3143.590 799.410 3144.770 ;
        RECT 796.630 3141.990 797.810 3143.170 ;
        RECT 798.230 3141.990 799.410 3143.170 ;
        RECT 796.630 2963.590 797.810 2964.770 ;
        RECT 798.230 2963.590 799.410 2964.770 ;
        RECT 796.630 2961.990 797.810 2963.170 ;
        RECT 798.230 2961.990 799.410 2963.170 ;
        RECT 796.630 2783.590 797.810 2784.770 ;
        RECT 798.230 2783.590 799.410 2784.770 ;
        RECT 796.630 2781.990 797.810 2783.170 ;
        RECT 798.230 2781.990 799.410 2783.170 ;
        RECT 796.630 2603.590 797.810 2604.770 ;
        RECT 798.230 2603.590 799.410 2604.770 ;
        RECT 796.630 2601.990 797.810 2603.170 ;
        RECT 798.230 2601.990 799.410 2603.170 ;
        RECT 796.630 2423.590 797.810 2424.770 ;
        RECT 798.230 2423.590 799.410 2424.770 ;
        RECT 796.630 2421.990 797.810 2423.170 ;
        RECT 798.230 2421.990 799.410 2423.170 ;
        RECT 796.630 2243.590 797.810 2244.770 ;
        RECT 798.230 2243.590 799.410 2244.770 ;
        RECT 796.630 2241.990 797.810 2243.170 ;
        RECT 798.230 2241.990 799.410 2243.170 ;
        RECT 796.630 2063.590 797.810 2064.770 ;
        RECT 798.230 2063.590 799.410 2064.770 ;
        RECT 796.630 2061.990 797.810 2063.170 ;
        RECT 798.230 2061.990 799.410 2063.170 ;
        RECT 796.630 1883.590 797.810 1884.770 ;
        RECT 798.230 1883.590 799.410 1884.770 ;
        RECT 796.630 1881.990 797.810 1883.170 ;
        RECT 798.230 1881.990 799.410 1883.170 ;
        RECT 796.630 1703.590 797.810 1704.770 ;
        RECT 798.230 1703.590 799.410 1704.770 ;
        RECT 796.630 1701.990 797.810 1703.170 ;
        RECT 798.230 1701.990 799.410 1703.170 ;
        RECT 796.630 1523.590 797.810 1524.770 ;
        RECT 798.230 1523.590 799.410 1524.770 ;
        RECT 796.630 1521.990 797.810 1523.170 ;
        RECT 798.230 1521.990 799.410 1523.170 ;
        RECT 796.630 1343.590 797.810 1344.770 ;
        RECT 798.230 1343.590 799.410 1344.770 ;
        RECT 796.630 1341.990 797.810 1343.170 ;
        RECT 798.230 1341.990 799.410 1343.170 ;
        RECT 796.630 1163.590 797.810 1164.770 ;
        RECT 798.230 1163.590 799.410 1164.770 ;
        RECT 796.630 1161.990 797.810 1163.170 ;
        RECT 798.230 1161.990 799.410 1163.170 ;
        RECT 796.630 983.590 797.810 984.770 ;
        RECT 798.230 983.590 799.410 984.770 ;
        RECT 796.630 981.990 797.810 983.170 ;
        RECT 798.230 981.990 799.410 983.170 ;
        RECT 796.630 803.590 797.810 804.770 ;
        RECT 798.230 803.590 799.410 804.770 ;
        RECT 796.630 801.990 797.810 803.170 ;
        RECT 798.230 801.990 799.410 803.170 ;
        RECT 256.630 623.590 257.810 624.770 ;
        RECT 258.230 623.590 259.410 624.770 ;
        RECT 256.630 621.990 257.810 623.170 ;
        RECT 258.230 621.990 259.410 623.170 ;
        RECT 796.630 623.590 797.810 624.770 ;
        RECT 798.230 623.590 799.410 624.770 ;
        RECT 796.630 621.990 797.810 623.170 ;
        RECT 798.230 621.990 799.410 623.170 ;
        RECT 256.630 443.590 257.810 444.770 ;
        RECT 258.230 443.590 259.410 444.770 ;
        RECT 256.630 441.990 257.810 443.170 ;
        RECT 258.230 441.990 259.410 443.170 ;
        RECT 256.630 263.590 257.810 264.770 ;
        RECT 258.230 263.590 259.410 264.770 ;
        RECT 256.630 261.990 257.810 263.170 ;
        RECT 258.230 261.990 259.410 263.170 ;
        RECT 256.630 83.590 257.810 84.770 ;
        RECT 258.230 83.590 259.410 84.770 ;
        RECT 256.630 81.990 257.810 83.170 ;
        RECT 258.230 81.990 259.410 83.170 ;
        RECT 256.630 -18.860 257.810 -17.680 ;
        RECT 258.230 -18.860 259.410 -17.680 ;
        RECT 256.630 -20.460 257.810 -19.280 ;
        RECT 258.230 -20.460 259.410 -19.280 ;
        RECT 436.630 443.590 437.810 444.770 ;
        RECT 438.230 443.590 439.410 444.770 ;
        RECT 436.630 441.990 437.810 443.170 ;
        RECT 438.230 441.990 439.410 443.170 ;
        RECT 436.630 263.590 437.810 264.770 ;
        RECT 438.230 263.590 439.410 264.770 ;
        RECT 436.630 261.990 437.810 263.170 ;
        RECT 438.230 261.990 439.410 263.170 ;
        RECT 436.630 83.590 437.810 84.770 ;
        RECT 438.230 83.590 439.410 84.770 ;
        RECT 436.630 81.990 437.810 83.170 ;
        RECT 438.230 81.990 439.410 83.170 ;
        RECT 436.630 -18.860 437.810 -17.680 ;
        RECT 438.230 -18.860 439.410 -17.680 ;
        RECT 436.630 -20.460 437.810 -19.280 ;
        RECT 438.230 -20.460 439.410 -19.280 ;
        RECT 616.630 443.590 617.810 444.770 ;
        RECT 618.230 443.590 619.410 444.770 ;
        RECT 616.630 441.990 617.810 443.170 ;
        RECT 618.230 441.990 619.410 443.170 ;
        RECT 616.630 263.590 617.810 264.770 ;
        RECT 618.230 263.590 619.410 264.770 ;
        RECT 616.630 261.990 617.810 263.170 ;
        RECT 618.230 261.990 619.410 263.170 ;
        RECT 616.630 83.590 617.810 84.770 ;
        RECT 618.230 83.590 619.410 84.770 ;
        RECT 616.630 81.990 617.810 83.170 ;
        RECT 618.230 81.990 619.410 83.170 ;
        RECT 616.630 -18.860 617.810 -17.680 ;
        RECT 618.230 -18.860 619.410 -17.680 ;
        RECT 616.630 -20.460 617.810 -19.280 ;
        RECT 618.230 -20.460 619.410 -19.280 ;
        RECT 796.630 443.590 797.810 444.770 ;
        RECT 798.230 443.590 799.410 444.770 ;
        RECT 796.630 441.990 797.810 443.170 ;
        RECT 798.230 441.990 799.410 443.170 ;
        RECT 796.630 263.590 797.810 264.770 ;
        RECT 798.230 263.590 799.410 264.770 ;
        RECT 796.630 261.990 797.810 263.170 ;
        RECT 798.230 261.990 799.410 263.170 ;
        RECT 796.630 83.590 797.810 84.770 ;
        RECT 798.230 83.590 799.410 84.770 ;
        RECT 796.630 81.990 797.810 83.170 ;
        RECT 798.230 81.990 799.410 83.170 ;
        RECT 796.630 -18.860 797.810 -17.680 ;
        RECT 798.230 -18.860 799.410 -17.680 ;
        RECT 796.630 -20.460 797.810 -19.280 ;
        RECT 798.230 -20.460 799.410 -19.280 ;
        RECT 976.630 3538.960 977.810 3540.140 ;
        RECT 978.230 3538.960 979.410 3540.140 ;
        RECT 976.630 3537.360 977.810 3538.540 ;
        RECT 978.230 3537.360 979.410 3538.540 ;
        RECT 976.630 3503.590 977.810 3504.770 ;
        RECT 978.230 3503.590 979.410 3504.770 ;
        RECT 976.630 3501.990 977.810 3503.170 ;
        RECT 978.230 3501.990 979.410 3503.170 ;
        RECT 976.630 3323.590 977.810 3324.770 ;
        RECT 978.230 3323.590 979.410 3324.770 ;
        RECT 976.630 3321.990 977.810 3323.170 ;
        RECT 978.230 3321.990 979.410 3323.170 ;
        RECT 976.630 3143.590 977.810 3144.770 ;
        RECT 978.230 3143.590 979.410 3144.770 ;
        RECT 976.630 3141.990 977.810 3143.170 ;
        RECT 978.230 3141.990 979.410 3143.170 ;
        RECT 976.630 2963.590 977.810 2964.770 ;
        RECT 978.230 2963.590 979.410 2964.770 ;
        RECT 976.630 2961.990 977.810 2963.170 ;
        RECT 978.230 2961.990 979.410 2963.170 ;
        RECT 976.630 2783.590 977.810 2784.770 ;
        RECT 978.230 2783.590 979.410 2784.770 ;
        RECT 976.630 2781.990 977.810 2783.170 ;
        RECT 978.230 2781.990 979.410 2783.170 ;
        RECT 976.630 2603.590 977.810 2604.770 ;
        RECT 978.230 2603.590 979.410 2604.770 ;
        RECT 976.630 2601.990 977.810 2603.170 ;
        RECT 978.230 2601.990 979.410 2603.170 ;
        RECT 976.630 2423.590 977.810 2424.770 ;
        RECT 978.230 2423.590 979.410 2424.770 ;
        RECT 976.630 2421.990 977.810 2423.170 ;
        RECT 978.230 2421.990 979.410 2423.170 ;
        RECT 976.630 2243.590 977.810 2244.770 ;
        RECT 978.230 2243.590 979.410 2244.770 ;
        RECT 976.630 2241.990 977.810 2243.170 ;
        RECT 978.230 2241.990 979.410 2243.170 ;
        RECT 976.630 2063.590 977.810 2064.770 ;
        RECT 978.230 2063.590 979.410 2064.770 ;
        RECT 976.630 2061.990 977.810 2063.170 ;
        RECT 978.230 2061.990 979.410 2063.170 ;
        RECT 976.630 1883.590 977.810 1884.770 ;
        RECT 978.230 1883.590 979.410 1884.770 ;
        RECT 976.630 1881.990 977.810 1883.170 ;
        RECT 978.230 1881.990 979.410 1883.170 ;
        RECT 976.630 1703.590 977.810 1704.770 ;
        RECT 978.230 1703.590 979.410 1704.770 ;
        RECT 976.630 1701.990 977.810 1703.170 ;
        RECT 978.230 1701.990 979.410 1703.170 ;
        RECT 976.630 1523.590 977.810 1524.770 ;
        RECT 978.230 1523.590 979.410 1524.770 ;
        RECT 976.630 1521.990 977.810 1523.170 ;
        RECT 978.230 1521.990 979.410 1523.170 ;
        RECT 976.630 1343.590 977.810 1344.770 ;
        RECT 978.230 1343.590 979.410 1344.770 ;
        RECT 976.630 1341.990 977.810 1343.170 ;
        RECT 978.230 1341.990 979.410 1343.170 ;
        RECT 976.630 1163.590 977.810 1164.770 ;
        RECT 978.230 1163.590 979.410 1164.770 ;
        RECT 976.630 1161.990 977.810 1163.170 ;
        RECT 978.230 1161.990 979.410 1163.170 ;
        RECT 976.630 983.590 977.810 984.770 ;
        RECT 978.230 983.590 979.410 984.770 ;
        RECT 976.630 981.990 977.810 983.170 ;
        RECT 978.230 981.990 979.410 983.170 ;
        RECT 976.630 803.590 977.810 804.770 ;
        RECT 978.230 803.590 979.410 804.770 ;
        RECT 976.630 801.990 977.810 803.170 ;
        RECT 978.230 801.990 979.410 803.170 ;
        RECT 976.630 623.590 977.810 624.770 ;
        RECT 978.230 623.590 979.410 624.770 ;
        RECT 976.630 621.990 977.810 623.170 ;
        RECT 978.230 621.990 979.410 623.170 ;
        RECT 976.630 443.590 977.810 444.770 ;
        RECT 978.230 443.590 979.410 444.770 ;
        RECT 976.630 441.990 977.810 443.170 ;
        RECT 978.230 441.990 979.410 443.170 ;
        RECT 976.630 263.590 977.810 264.770 ;
        RECT 978.230 263.590 979.410 264.770 ;
        RECT 976.630 261.990 977.810 263.170 ;
        RECT 978.230 261.990 979.410 263.170 ;
        RECT 976.630 83.590 977.810 84.770 ;
        RECT 978.230 83.590 979.410 84.770 ;
        RECT 976.630 81.990 977.810 83.170 ;
        RECT 978.230 81.990 979.410 83.170 ;
        RECT 976.630 -18.860 977.810 -17.680 ;
        RECT 978.230 -18.860 979.410 -17.680 ;
        RECT 976.630 -20.460 977.810 -19.280 ;
        RECT 978.230 -20.460 979.410 -19.280 ;
        RECT 1156.630 3538.960 1157.810 3540.140 ;
        RECT 1158.230 3538.960 1159.410 3540.140 ;
        RECT 1156.630 3537.360 1157.810 3538.540 ;
        RECT 1158.230 3537.360 1159.410 3538.540 ;
        RECT 1156.630 3503.590 1157.810 3504.770 ;
        RECT 1158.230 3503.590 1159.410 3504.770 ;
        RECT 1156.630 3501.990 1157.810 3503.170 ;
        RECT 1158.230 3501.990 1159.410 3503.170 ;
        RECT 1156.630 3323.590 1157.810 3324.770 ;
        RECT 1158.230 3323.590 1159.410 3324.770 ;
        RECT 1156.630 3321.990 1157.810 3323.170 ;
        RECT 1158.230 3321.990 1159.410 3323.170 ;
        RECT 1156.630 3143.590 1157.810 3144.770 ;
        RECT 1158.230 3143.590 1159.410 3144.770 ;
        RECT 1156.630 3141.990 1157.810 3143.170 ;
        RECT 1158.230 3141.990 1159.410 3143.170 ;
        RECT 1156.630 2963.590 1157.810 2964.770 ;
        RECT 1158.230 2963.590 1159.410 2964.770 ;
        RECT 1156.630 2961.990 1157.810 2963.170 ;
        RECT 1158.230 2961.990 1159.410 2963.170 ;
        RECT 1156.630 2783.590 1157.810 2784.770 ;
        RECT 1158.230 2783.590 1159.410 2784.770 ;
        RECT 1156.630 2781.990 1157.810 2783.170 ;
        RECT 1158.230 2781.990 1159.410 2783.170 ;
        RECT 1156.630 2603.590 1157.810 2604.770 ;
        RECT 1158.230 2603.590 1159.410 2604.770 ;
        RECT 1156.630 2601.990 1157.810 2603.170 ;
        RECT 1158.230 2601.990 1159.410 2603.170 ;
        RECT 1156.630 2423.590 1157.810 2424.770 ;
        RECT 1158.230 2423.590 1159.410 2424.770 ;
        RECT 1156.630 2421.990 1157.810 2423.170 ;
        RECT 1158.230 2421.990 1159.410 2423.170 ;
        RECT 1156.630 2243.590 1157.810 2244.770 ;
        RECT 1158.230 2243.590 1159.410 2244.770 ;
        RECT 1156.630 2241.990 1157.810 2243.170 ;
        RECT 1158.230 2241.990 1159.410 2243.170 ;
        RECT 1156.630 2063.590 1157.810 2064.770 ;
        RECT 1158.230 2063.590 1159.410 2064.770 ;
        RECT 1156.630 2061.990 1157.810 2063.170 ;
        RECT 1158.230 2061.990 1159.410 2063.170 ;
        RECT 1156.630 1883.590 1157.810 1884.770 ;
        RECT 1158.230 1883.590 1159.410 1884.770 ;
        RECT 1156.630 1881.990 1157.810 1883.170 ;
        RECT 1158.230 1881.990 1159.410 1883.170 ;
        RECT 1156.630 1703.590 1157.810 1704.770 ;
        RECT 1158.230 1703.590 1159.410 1704.770 ;
        RECT 1156.630 1701.990 1157.810 1703.170 ;
        RECT 1158.230 1701.990 1159.410 1703.170 ;
        RECT 1156.630 1523.590 1157.810 1524.770 ;
        RECT 1158.230 1523.590 1159.410 1524.770 ;
        RECT 1156.630 1521.990 1157.810 1523.170 ;
        RECT 1158.230 1521.990 1159.410 1523.170 ;
        RECT 1156.630 1343.590 1157.810 1344.770 ;
        RECT 1158.230 1343.590 1159.410 1344.770 ;
        RECT 1156.630 1341.990 1157.810 1343.170 ;
        RECT 1158.230 1341.990 1159.410 1343.170 ;
        RECT 1156.630 1163.590 1157.810 1164.770 ;
        RECT 1158.230 1163.590 1159.410 1164.770 ;
        RECT 1156.630 1161.990 1157.810 1163.170 ;
        RECT 1158.230 1161.990 1159.410 1163.170 ;
        RECT 1156.630 983.590 1157.810 984.770 ;
        RECT 1158.230 983.590 1159.410 984.770 ;
        RECT 1156.630 981.990 1157.810 983.170 ;
        RECT 1158.230 981.990 1159.410 983.170 ;
        RECT 1156.630 803.590 1157.810 804.770 ;
        RECT 1158.230 803.590 1159.410 804.770 ;
        RECT 1156.630 801.990 1157.810 803.170 ;
        RECT 1158.230 801.990 1159.410 803.170 ;
        RECT 1156.630 623.590 1157.810 624.770 ;
        RECT 1158.230 623.590 1159.410 624.770 ;
        RECT 1156.630 621.990 1157.810 623.170 ;
        RECT 1158.230 621.990 1159.410 623.170 ;
        RECT 1156.630 443.590 1157.810 444.770 ;
        RECT 1158.230 443.590 1159.410 444.770 ;
        RECT 1156.630 441.990 1157.810 443.170 ;
        RECT 1158.230 441.990 1159.410 443.170 ;
        RECT 1156.630 263.590 1157.810 264.770 ;
        RECT 1158.230 263.590 1159.410 264.770 ;
        RECT 1156.630 261.990 1157.810 263.170 ;
        RECT 1158.230 261.990 1159.410 263.170 ;
        RECT 1156.630 83.590 1157.810 84.770 ;
        RECT 1158.230 83.590 1159.410 84.770 ;
        RECT 1156.630 81.990 1157.810 83.170 ;
        RECT 1158.230 81.990 1159.410 83.170 ;
        RECT 1156.630 -18.860 1157.810 -17.680 ;
        RECT 1158.230 -18.860 1159.410 -17.680 ;
        RECT 1156.630 -20.460 1157.810 -19.280 ;
        RECT 1158.230 -20.460 1159.410 -19.280 ;
        RECT 1336.630 3538.960 1337.810 3540.140 ;
        RECT 1338.230 3538.960 1339.410 3540.140 ;
        RECT 1336.630 3537.360 1337.810 3538.540 ;
        RECT 1338.230 3537.360 1339.410 3538.540 ;
        RECT 1336.630 3503.590 1337.810 3504.770 ;
        RECT 1338.230 3503.590 1339.410 3504.770 ;
        RECT 1336.630 3501.990 1337.810 3503.170 ;
        RECT 1338.230 3501.990 1339.410 3503.170 ;
        RECT 1336.630 3323.590 1337.810 3324.770 ;
        RECT 1338.230 3323.590 1339.410 3324.770 ;
        RECT 1336.630 3321.990 1337.810 3323.170 ;
        RECT 1338.230 3321.990 1339.410 3323.170 ;
        RECT 1336.630 3143.590 1337.810 3144.770 ;
        RECT 1338.230 3143.590 1339.410 3144.770 ;
        RECT 1336.630 3141.990 1337.810 3143.170 ;
        RECT 1338.230 3141.990 1339.410 3143.170 ;
        RECT 1336.630 2963.590 1337.810 2964.770 ;
        RECT 1338.230 2963.590 1339.410 2964.770 ;
        RECT 1336.630 2961.990 1337.810 2963.170 ;
        RECT 1338.230 2961.990 1339.410 2963.170 ;
        RECT 1336.630 2783.590 1337.810 2784.770 ;
        RECT 1338.230 2783.590 1339.410 2784.770 ;
        RECT 1336.630 2781.990 1337.810 2783.170 ;
        RECT 1338.230 2781.990 1339.410 2783.170 ;
        RECT 1336.630 2603.590 1337.810 2604.770 ;
        RECT 1338.230 2603.590 1339.410 2604.770 ;
        RECT 1336.630 2601.990 1337.810 2603.170 ;
        RECT 1338.230 2601.990 1339.410 2603.170 ;
        RECT 1336.630 2423.590 1337.810 2424.770 ;
        RECT 1338.230 2423.590 1339.410 2424.770 ;
        RECT 1336.630 2421.990 1337.810 2423.170 ;
        RECT 1338.230 2421.990 1339.410 2423.170 ;
        RECT 1336.630 2243.590 1337.810 2244.770 ;
        RECT 1338.230 2243.590 1339.410 2244.770 ;
        RECT 1336.630 2241.990 1337.810 2243.170 ;
        RECT 1338.230 2241.990 1339.410 2243.170 ;
        RECT 1336.630 2063.590 1337.810 2064.770 ;
        RECT 1338.230 2063.590 1339.410 2064.770 ;
        RECT 1336.630 2061.990 1337.810 2063.170 ;
        RECT 1338.230 2061.990 1339.410 2063.170 ;
        RECT 1336.630 1883.590 1337.810 1884.770 ;
        RECT 1338.230 1883.590 1339.410 1884.770 ;
        RECT 1336.630 1881.990 1337.810 1883.170 ;
        RECT 1338.230 1881.990 1339.410 1883.170 ;
        RECT 1336.630 1703.590 1337.810 1704.770 ;
        RECT 1338.230 1703.590 1339.410 1704.770 ;
        RECT 1336.630 1701.990 1337.810 1703.170 ;
        RECT 1338.230 1701.990 1339.410 1703.170 ;
        RECT 1336.630 1523.590 1337.810 1524.770 ;
        RECT 1338.230 1523.590 1339.410 1524.770 ;
        RECT 1336.630 1521.990 1337.810 1523.170 ;
        RECT 1338.230 1521.990 1339.410 1523.170 ;
        RECT 1336.630 1343.590 1337.810 1344.770 ;
        RECT 1338.230 1343.590 1339.410 1344.770 ;
        RECT 1336.630 1341.990 1337.810 1343.170 ;
        RECT 1338.230 1341.990 1339.410 1343.170 ;
        RECT 1336.630 1163.590 1337.810 1164.770 ;
        RECT 1338.230 1163.590 1339.410 1164.770 ;
        RECT 1336.630 1161.990 1337.810 1163.170 ;
        RECT 1338.230 1161.990 1339.410 1163.170 ;
        RECT 1336.630 983.590 1337.810 984.770 ;
        RECT 1338.230 983.590 1339.410 984.770 ;
        RECT 1336.630 981.990 1337.810 983.170 ;
        RECT 1338.230 981.990 1339.410 983.170 ;
        RECT 1336.630 803.590 1337.810 804.770 ;
        RECT 1338.230 803.590 1339.410 804.770 ;
        RECT 1336.630 801.990 1337.810 803.170 ;
        RECT 1338.230 801.990 1339.410 803.170 ;
        RECT 1336.630 623.590 1337.810 624.770 ;
        RECT 1338.230 623.590 1339.410 624.770 ;
        RECT 1336.630 621.990 1337.810 623.170 ;
        RECT 1338.230 621.990 1339.410 623.170 ;
        RECT 1336.630 443.590 1337.810 444.770 ;
        RECT 1338.230 443.590 1339.410 444.770 ;
        RECT 1336.630 441.990 1337.810 443.170 ;
        RECT 1338.230 441.990 1339.410 443.170 ;
        RECT 1336.630 263.590 1337.810 264.770 ;
        RECT 1338.230 263.590 1339.410 264.770 ;
        RECT 1336.630 261.990 1337.810 263.170 ;
        RECT 1338.230 261.990 1339.410 263.170 ;
        RECT 1336.630 83.590 1337.810 84.770 ;
        RECT 1338.230 83.590 1339.410 84.770 ;
        RECT 1336.630 81.990 1337.810 83.170 ;
        RECT 1338.230 81.990 1339.410 83.170 ;
        RECT 1336.630 -18.860 1337.810 -17.680 ;
        RECT 1338.230 -18.860 1339.410 -17.680 ;
        RECT 1336.630 -20.460 1337.810 -19.280 ;
        RECT 1338.230 -20.460 1339.410 -19.280 ;
        RECT 1516.630 3538.960 1517.810 3540.140 ;
        RECT 1518.230 3538.960 1519.410 3540.140 ;
        RECT 1516.630 3537.360 1517.810 3538.540 ;
        RECT 1518.230 3537.360 1519.410 3538.540 ;
        RECT 1516.630 3503.590 1517.810 3504.770 ;
        RECT 1518.230 3503.590 1519.410 3504.770 ;
        RECT 1516.630 3501.990 1517.810 3503.170 ;
        RECT 1518.230 3501.990 1519.410 3503.170 ;
        RECT 1516.630 3323.590 1517.810 3324.770 ;
        RECT 1518.230 3323.590 1519.410 3324.770 ;
        RECT 1516.630 3321.990 1517.810 3323.170 ;
        RECT 1518.230 3321.990 1519.410 3323.170 ;
        RECT 1516.630 3143.590 1517.810 3144.770 ;
        RECT 1518.230 3143.590 1519.410 3144.770 ;
        RECT 1516.630 3141.990 1517.810 3143.170 ;
        RECT 1518.230 3141.990 1519.410 3143.170 ;
        RECT 1516.630 2963.590 1517.810 2964.770 ;
        RECT 1518.230 2963.590 1519.410 2964.770 ;
        RECT 1516.630 2961.990 1517.810 2963.170 ;
        RECT 1518.230 2961.990 1519.410 2963.170 ;
        RECT 1516.630 2783.590 1517.810 2784.770 ;
        RECT 1518.230 2783.590 1519.410 2784.770 ;
        RECT 1516.630 2781.990 1517.810 2783.170 ;
        RECT 1518.230 2781.990 1519.410 2783.170 ;
        RECT 1516.630 2603.590 1517.810 2604.770 ;
        RECT 1518.230 2603.590 1519.410 2604.770 ;
        RECT 1516.630 2601.990 1517.810 2603.170 ;
        RECT 1518.230 2601.990 1519.410 2603.170 ;
        RECT 1516.630 2423.590 1517.810 2424.770 ;
        RECT 1518.230 2423.590 1519.410 2424.770 ;
        RECT 1516.630 2421.990 1517.810 2423.170 ;
        RECT 1518.230 2421.990 1519.410 2423.170 ;
        RECT 1516.630 2243.590 1517.810 2244.770 ;
        RECT 1518.230 2243.590 1519.410 2244.770 ;
        RECT 1516.630 2241.990 1517.810 2243.170 ;
        RECT 1518.230 2241.990 1519.410 2243.170 ;
        RECT 1516.630 2063.590 1517.810 2064.770 ;
        RECT 1518.230 2063.590 1519.410 2064.770 ;
        RECT 1516.630 2061.990 1517.810 2063.170 ;
        RECT 1518.230 2061.990 1519.410 2063.170 ;
        RECT 1516.630 1883.590 1517.810 1884.770 ;
        RECT 1518.230 1883.590 1519.410 1884.770 ;
        RECT 1516.630 1881.990 1517.810 1883.170 ;
        RECT 1518.230 1881.990 1519.410 1883.170 ;
        RECT 1516.630 1703.590 1517.810 1704.770 ;
        RECT 1518.230 1703.590 1519.410 1704.770 ;
        RECT 1516.630 1701.990 1517.810 1703.170 ;
        RECT 1518.230 1701.990 1519.410 1703.170 ;
        RECT 1516.630 1523.590 1517.810 1524.770 ;
        RECT 1518.230 1523.590 1519.410 1524.770 ;
        RECT 1516.630 1521.990 1517.810 1523.170 ;
        RECT 1518.230 1521.990 1519.410 1523.170 ;
        RECT 1516.630 1343.590 1517.810 1344.770 ;
        RECT 1518.230 1343.590 1519.410 1344.770 ;
        RECT 1516.630 1341.990 1517.810 1343.170 ;
        RECT 1518.230 1341.990 1519.410 1343.170 ;
        RECT 1516.630 1163.590 1517.810 1164.770 ;
        RECT 1518.230 1163.590 1519.410 1164.770 ;
        RECT 1516.630 1161.990 1517.810 1163.170 ;
        RECT 1518.230 1161.990 1519.410 1163.170 ;
        RECT 1516.630 983.590 1517.810 984.770 ;
        RECT 1518.230 983.590 1519.410 984.770 ;
        RECT 1516.630 981.990 1517.810 983.170 ;
        RECT 1518.230 981.990 1519.410 983.170 ;
        RECT 1516.630 803.590 1517.810 804.770 ;
        RECT 1518.230 803.590 1519.410 804.770 ;
        RECT 1516.630 801.990 1517.810 803.170 ;
        RECT 1518.230 801.990 1519.410 803.170 ;
        RECT 1516.630 623.590 1517.810 624.770 ;
        RECT 1518.230 623.590 1519.410 624.770 ;
        RECT 1516.630 621.990 1517.810 623.170 ;
        RECT 1518.230 621.990 1519.410 623.170 ;
        RECT 1516.630 443.590 1517.810 444.770 ;
        RECT 1518.230 443.590 1519.410 444.770 ;
        RECT 1516.630 441.990 1517.810 443.170 ;
        RECT 1518.230 441.990 1519.410 443.170 ;
        RECT 1516.630 263.590 1517.810 264.770 ;
        RECT 1518.230 263.590 1519.410 264.770 ;
        RECT 1516.630 261.990 1517.810 263.170 ;
        RECT 1518.230 261.990 1519.410 263.170 ;
        RECT 1516.630 83.590 1517.810 84.770 ;
        RECT 1518.230 83.590 1519.410 84.770 ;
        RECT 1516.630 81.990 1517.810 83.170 ;
        RECT 1518.230 81.990 1519.410 83.170 ;
        RECT 1516.630 -18.860 1517.810 -17.680 ;
        RECT 1518.230 -18.860 1519.410 -17.680 ;
        RECT 1516.630 -20.460 1517.810 -19.280 ;
        RECT 1518.230 -20.460 1519.410 -19.280 ;
        RECT 1696.630 3538.960 1697.810 3540.140 ;
        RECT 1698.230 3538.960 1699.410 3540.140 ;
        RECT 1696.630 3537.360 1697.810 3538.540 ;
        RECT 1698.230 3537.360 1699.410 3538.540 ;
        RECT 1696.630 3503.590 1697.810 3504.770 ;
        RECT 1698.230 3503.590 1699.410 3504.770 ;
        RECT 1696.630 3501.990 1697.810 3503.170 ;
        RECT 1698.230 3501.990 1699.410 3503.170 ;
        RECT 1696.630 3323.590 1697.810 3324.770 ;
        RECT 1698.230 3323.590 1699.410 3324.770 ;
        RECT 1696.630 3321.990 1697.810 3323.170 ;
        RECT 1698.230 3321.990 1699.410 3323.170 ;
        RECT 1696.630 3143.590 1697.810 3144.770 ;
        RECT 1698.230 3143.590 1699.410 3144.770 ;
        RECT 1696.630 3141.990 1697.810 3143.170 ;
        RECT 1698.230 3141.990 1699.410 3143.170 ;
        RECT 1696.630 2963.590 1697.810 2964.770 ;
        RECT 1698.230 2963.590 1699.410 2964.770 ;
        RECT 1696.630 2961.990 1697.810 2963.170 ;
        RECT 1698.230 2961.990 1699.410 2963.170 ;
        RECT 1696.630 2783.590 1697.810 2784.770 ;
        RECT 1698.230 2783.590 1699.410 2784.770 ;
        RECT 1696.630 2781.990 1697.810 2783.170 ;
        RECT 1698.230 2781.990 1699.410 2783.170 ;
        RECT 1696.630 2603.590 1697.810 2604.770 ;
        RECT 1698.230 2603.590 1699.410 2604.770 ;
        RECT 1696.630 2601.990 1697.810 2603.170 ;
        RECT 1698.230 2601.990 1699.410 2603.170 ;
        RECT 1696.630 2423.590 1697.810 2424.770 ;
        RECT 1698.230 2423.590 1699.410 2424.770 ;
        RECT 1696.630 2421.990 1697.810 2423.170 ;
        RECT 1698.230 2421.990 1699.410 2423.170 ;
        RECT 1696.630 2243.590 1697.810 2244.770 ;
        RECT 1698.230 2243.590 1699.410 2244.770 ;
        RECT 1696.630 2241.990 1697.810 2243.170 ;
        RECT 1698.230 2241.990 1699.410 2243.170 ;
        RECT 1696.630 2063.590 1697.810 2064.770 ;
        RECT 1698.230 2063.590 1699.410 2064.770 ;
        RECT 1696.630 2061.990 1697.810 2063.170 ;
        RECT 1698.230 2061.990 1699.410 2063.170 ;
        RECT 1696.630 1883.590 1697.810 1884.770 ;
        RECT 1698.230 1883.590 1699.410 1884.770 ;
        RECT 1696.630 1881.990 1697.810 1883.170 ;
        RECT 1698.230 1881.990 1699.410 1883.170 ;
        RECT 1696.630 1703.590 1697.810 1704.770 ;
        RECT 1698.230 1703.590 1699.410 1704.770 ;
        RECT 1696.630 1701.990 1697.810 1703.170 ;
        RECT 1698.230 1701.990 1699.410 1703.170 ;
        RECT 1696.630 1523.590 1697.810 1524.770 ;
        RECT 1698.230 1523.590 1699.410 1524.770 ;
        RECT 1696.630 1521.990 1697.810 1523.170 ;
        RECT 1698.230 1521.990 1699.410 1523.170 ;
        RECT 1696.630 1343.590 1697.810 1344.770 ;
        RECT 1698.230 1343.590 1699.410 1344.770 ;
        RECT 1696.630 1341.990 1697.810 1343.170 ;
        RECT 1698.230 1341.990 1699.410 1343.170 ;
        RECT 1696.630 1163.590 1697.810 1164.770 ;
        RECT 1698.230 1163.590 1699.410 1164.770 ;
        RECT 1696.630 1161.990 1697.810 1163.170 ;
        RECT 1698.230 1161.990 1699.410 1163.170 ;
        RECT 1696.630 983.590 1697.810 984.770 ;
        RECT 1698.230 983.590 1699.410 984.770 ;
        RECT 1696.630 981.990 1697.810 983.170 ;
        RECT 1698.230 981.990 1699.410 983.170 ;
        RECT 1696.630 803.590 1697.810 804.770 ;
        RECT 1698.230 803.590 1699.410 804.770 ;
        RECT 1696.630 801.990 1697.810 803.170 ;
        RECT 1698.230 801.990 1699.410 803.170 ;
        RECT 1696.630 623.590 1697.810 624.770 ;
        RECT 1698.230 623.590 1699.410 624.770 ;
        RECT 1696.630 621.990 1697.810 623.170 ;
        RECT 1698.230 621.990 1699.410 623.170 ;
        RECT 1696.630 443.590 1697.810 444.770 ;
        RECT 1698.230 443.590 1699.410 444.770 ;
        RECT 1696.630 441.990 1697.810 443.170 ;
        RECT 1698.230 441.990 1699.410 443.170 ;
        RECT 1696.630 263.590 1697.810 264.770 ;
        RECT 1698.230 263.590 1699.410 264.770 ;
        RECT 1696.630 261.990 1697.810 263.170 ;
        RECT 1698.230 261.990 1699.410 263.170 ;
        RECT 1696.630 83.590 1697.810 84.770 ;
        RECT 1698.230 83.590 1699.410 84.770 ;
        RECT 1696.630 81.990 1697.810 83.170 ;
        RECT 1698.230 81.990 1699.410 83.170 ;
        RECT 1696.630 -18.860 1697.810 -17.680 ;
        RECT 1698.230 -18.860 1699.410 -17.680 ;
        RECT 1696.630 -20.460 1697.810 -19.280 ;
        RECT 1698.230 -20.460 1699.410 -19.280 ;
        RECT 1876.630 3538.960 1877.810 3540.140 ;
        RECT 1878.230 3538.960 1879.410 3540.140 ;
        RECT 1876.630 3537.360 1877.810 3538.540 ;
        RECT 1878.230 3537.360 1879.410 3538.540 ;
        RECT 1876.630 3503.590 1877.810 3504.770 ;
        RECT 1878.230 3503.590 1879.410 3504.770 ;
        RECT 1876.630 3501.990 1877.810 3503.170 ;
        RECT 1878.230 3501.990 1879.410 3503.170 ;
        RECT 1876.630 3323.590 1877.810 3324.770 ;
        RECT 1878.230 3323.590 1879.410 3324.770 ;
        RECT 1876.630 3321.990 1877.810 3323.170 ;
        RECT 1878.230 3321.990 1879.410 3323.170 ;
        RECT 1876.630 3143.590 1877.810 3144.770 ;
        RECT 1878.230 3143.590 1879.410 3144.770 ;
        RECT 1876.630 3141.990 1877.810 3143.170 ;
        RECT 1878.230 3141.990 1879.410 3143.170 ;
        RECT 1876.630 2963.590 1877.810 2964.770 ;
        RECT 1878.230 2963.590 1879.410 2964.770 ;
        RECT 1876.630 2961.990 1877.810 2963.170 ;
        RECT 1878.230 2961.990 1879.410 2963.170 ;
        RECT 1876.630 2783.590 1877.810 2784.770 ;
        RECT 1878.230 2783.590 1879.410 2784.770 ;
        RECT 1876.630 2781.990 1877.810 2783.170 ;
        RECT 1878.230 2781.990 1879.410 2783.170 ;
        RECT 1876.630 2603.590 1877.810 2604.770 ;
        RECT 1878.230 2603.590 1879.410 2604.770 ;
        RECT 1876.630 2601.990 1877.810 2603.170 ;
        RECT 1878.230 2601.990 1879.410 2603.170 ;
        RECT 1876.630 2423.590 1877.810 2424.770 ;
        RECT 1878.230 2423.590 1879.410 2424.770 ;
        RECT 1876.630 2421.990 1877.810 2423.170 ;
        RECT 1878.230 2421.990 1879.410 2423.170 ;
        RECT 1876.630 2243.590 1877.810 2244.770 ;
        RECT 1878.230 2243.590 1879.410 2244.770 ;
        RECT 1876.630 2241.990 1877.810 2243.170 ;
        RECT 1878.230 2241.990 1879.410 2243.170 ;
        RECT 1876.630 2063.590 1877.810 2064.770 ;
        RECT 1878.230 2063.590 1879.410 2064.770 ;
        RECT 1876.630 2061.990 1877.810 2063.170 ;
        RECT 1878.230 2061.990 1879.410 2063.170 ;
        RECT 1876.630 1883.590 1877.810 1884.770 ;
        RECT 1878.230 1883.590 1879.410 1884.770 ;
        RECT 1876.630 1881.990 1877.810 1883.170 ;
        RECT 1878.230 1881.990 1879.410 1883.170 ;
        RECT 1876.630 1703.590 1877.810 1704.770 ;
        RECT 1878.230 1703.590 1879.410 1704.770 ;
        RECT 1876.630 1701.990 1877.810 1703.170 ;
        RECT 1878.230 1701.990 1879.410 1703.170 ;
        RECT 1876.630 1523.590 1877.810 1524.770 ;
        RECT 1878.230 1523.590 1879.410 1524.770 ;
        RECT 1876.630 1521.990 1877.810 1523.170 ;
        RECT 1878.230 1521.990 1879.410 1523.170 ;
        RECT 1876.630 1343.590 1877.810 1344.770 ;
        RECT 1878.230 1343.590 1879.410 1344.770 ;
        RECT 1876.630 1341.990 1877.810 1343.170 ;
        RECT 1878.230 1341.990 1879.410 1343.170 ;
        RECT 1876.630 1163.590 1877.810 1164.770 ;
        RECT 1878.230 1163.590 1879.410 1164.770 ;
        RECT 1876.630 1161.990 1877.810 1163.170 ;
        RECT 1878.230 1161.990 1879.410 1163.170 ;
        RECT 1876.630 983.590 1877.810 984.770 ;
        RECT 1878.230 983.590 1879.410 984.770 ;
        RECT 1876.630 981.990 1877.810 983.170 ;
        RECT 1878.230 981.990 1879.410 983.170 ;
        RECT 1876.630 803.590 1877.810 804.770 ;
        RECT 1878.230 803.590 1879.410 804.770 ;
        RECT 1876.630 801.990 1877.810 803.170 ;
        RECT 1878.230 801.990 1879.410 803.170 ;
        RECT 1876.630 623.590 1877.810 624.770 ;
        RECT 1878.230 623.590 1879.410 624.770 ;
        RECT 1876.630 621.990 1877.810 623.170 ;
        RECT 1878.230 621.990 1879.410 623.170 ;
        RECT 1876.630 443.590 1877.810 444.770 ;
        RECT 1878.230 443.590 1879.410 444.770 ;
        RECT 1876.630 441.990 1877.810 443.170 ;
        RECT 1878.230 441.990 1879.410 443.170 ;
        RECT 1876.630 263.590 1877.810 264.770 ;
        RECT 1878.230 263.590 1879.410 264.770 ;
        RECT 1876.630 261.990 1877.810 263.170 ;
        RECT 1878.230 261.990 1879.410 263.170 ;
        RECT 1876.630 83.590 1877.810 84.770 ;
        RECT 1878.230 83.590 1879.410 84.770 ;
        RECT 1876.630 81.990 1877.810 83.170 ;
        RECT 1878.230 81.990 1879.410 83.170 ;
        RECT 1876.630 -18.860 1877.810 -17.680 ;
        RECT 1878.230 -18.860 1879.410 -17.680 ;
        RECT 1876.630 -20.460 1877.810 -19.280 ;
        RECT 1878.230 -20.460 1879.410 -19.280 ;
        RECT 2056.630 3538.960 2057.810 3540.140 ;
        RECT 2058.230 3538.960 2059.410 3540.140 ;
        RECT 2056.630 3537.360 2057.810 3538.540 ;
        RECT 2058.230 3537.360 2059.410 3538.540 ;
        RECT 2056.630 3503.590 2057.810 3504.770 ;
        RECT 2058.230 3503.590 2059.410 3504.770 ;
        RECT 2056.630 3501.990 2057.810 3503.170 ;
        RECT 2058.230 3501.990 2059.410 3503.170 ;
        RECT 2056.630 3323.590 2057.810 3324.770 ;
        RECT 2058.230 3323.590 2059.410 3324.770 ;
        RECT 2056.630 3321.990 2057.810 3323.170 ;
        RECT 2058.230 3321.990 2059.410 3323.170 ;
        RECT 2056.630 3143.590 2057.810 3144.770 ;
        RECT 2058.230 3143.590 2059.410 3144.770 ;
        RECT 2056.630 3141.990 2057.810 3143.170 ;
        RECT 2058.230 3141.990 2059.410 3143.170 ;
        RECT 2056.630 2963.590 2057.810 2964.770 ;
        RECT 2058.230 2963.590 2059.410 2964.770 ;
        RECT 2056.630 2961.990 2057.810 2963.170 ;
        RECT 2058.230 2961.990 2059.410 2963.170 ;
        RECT 2056.630 2783.590 2057.810 2784.770 ;
        RECT 2058.230 2783.590 2059.410 2784.770 ;
        RECT 2056.630 2781.990 2057.810 2783.170 ;
        RECT 2058.230 2781.990 2059.410 2783.170 ;
        RECT 2056.630 2603.590 2057.810 2604.770 ;
        RECT 2058.230 2603.590 2059.410 2604.770 ;
        RECT 2056.630 2601.990 2057.810 2603.170 ;
        RECT 2058.230 2601.990 2059.410 2603.170 ;
        RECT 2056.630 2423.590 2057.810 2424.770 ;
        RECT 2058.230 2423.590 2059.410 2424.770 ;
        RECT 2056.630 2421.990 2057.810 2423.170 ;
        RECT 2058.230 2421.990 2059.410 2423.170 ;
        RECT 2056.630 2243.590 2057.810 2244.770 ;
        RECT 2058.230 2243.590 2059.410 2244.770 ;
        RECT 2056.630 2241.990 2057.810 2243.170 ;
        RECT 2058.230 2241.990 2059.410 2243.170 ;
        RECT 2056.630 2063.590 2057.810 2064.770 ;
        RECT 2058.230 2063.590 2059.410 2064.770 ;
        RECT 2056.630 2061.990 2057.810 2063.170 ;
        RECT 2058.230 2061.990 2059.410 2063.170 ;
        RECT 2056.630 1883.590 2057.810 1884.770 ;
        RECT 2058.230 1883.590 2059.410 1884.770 ;
        RECT 2056.630 1881.990 2057.810 1883.170 ;
        RECT 2058.230 1881.990 2059.410 1883.170 ;
        RECT 2056.630 1703.590 2057.810 1704.770 ;
        RECT 2058.230 1703.590 2059.410 1704.770 ;
        RECT 2056.630 1701.990 2057.810 1703.170 ;
        RECT 2058.230 1701.990 2059.410 1703.170 ;
        RECT 2056.630 1523.590 2057.810 1524.770 ;
        RECT 2058.230 1523.590 2059.410 1524.770 ;
        RECT 2056.630 1521.990 2057.810 1523.170 ;
        RECT 2058.230 1521.990 2059.410 1523.170 ;
        RECT 2056.630 1343.590 2057.810 1344.770 ;
        RECT 2058.230 1343.590 2059.410 1344.770 ;
        RECT 2056.630 1341.990 2057.810 1343.170 ;
        RECT 2058.230 1341.990 2059.410 1343.170 ;
        RECT 2056.630 1163.590 2057.810 1164.770 ;
        RECT 2058.230 1163.590 2059.410 1164.770 ;
        RECT 2056.630 1161.990 2057.810 1163.170 ;
        RECT 2058.230 1161.990 2059.410 1163.170 ;
        RECT 2056.630 983.590 2057.810 984.770 ;
        RECT 2058.230 983.590 2059.410 984.770 ;
        RECT 2056.630 981.990 2057.810 983.170 ;
        RECT 2058.230 981.990 2059.410 983.170 ;
        RECT 2056.630 803.590 2057.810 804.770 ;
        RECT 2058.230 803.590 2059.410 804.770 ;
        RECT 2056.630 801.990 2057.810 803.170 ;
        RECT 2058.230 801.990 2059.410 803.170 ;
        RECT 2056.630 623.590 2057.810 624.770 ;
        RECT 2058.230 623.590 2059.410 624.770 ;
        RECT 2056.630 621.990 2057.810 623.170 ;
        RECT 2058.230 621.990 2059.410 623.170 ;
        RECT 2056.630 443.590 2057.810 444.770 ;
        RECT 2058.230 443.590 2059.410 444.770 ;
        RECT 2056.630 441.990 2057.810 443.170 ;
        RECT 2058.230 441.990 2059.410 443.170 ;
        RECT 2056.630 263.590 2057.810 264.770 ;
        RECT 2058.230 263.590 2059.410 264.770 ;
        RECT 2056.630 261.990 2057.810 263.170 ;
        RECT 2058.230 261.990 2059.410 263.170 ;
        RECT 2056.630 83.590 2057.810 84.770 ;
        RECT 2058.230 83.590 2059.410 84.770 ;
        RECT 2056.630 81.990 2057.810 83.170 ;
        RECT 2058.230 81.990 2059.410 83.170 ;
        RECT 2056.630 -18.860 2057.810 -17.680 ;
        RECT 2058.230 -18.860 2059.410 -17.680 ;
        RECT 2056.630 -20.460 2057.810 -19.280 ;
        RECT 2058.230 -20.460 2059.410 -19.280 ;
        RECT 2236.630 3538.960 2237.810 3540.140 ;
        RECT 2238.230 3538.960 2239.410 3540.140 ;
        RECT 2236.630 3537.360 2237.810 3538.540 ;
        RECT 2238.230 3537.360 2239.410 3538.540 ;
        RECT 2236.630 3503.590 2237.810 3504.770 ;
        RECT 2238.230 3503.590 2239.410 3504.770 ;
        RECT 2236.630 3501.990 2237.810 3503.170 ;
        RECT 2238.230 3501.990 2239.410 3503.170 ;
        RECT 2236.630 3323.590 2237.810 3324.770 ;
        RECT 2238.230 3323.590 2239.410 3324.770 ;
        RECT 2236.630 3321.990 2237.810 3323.170 ;
        RECT 2238.230 3321.990 2239.410 3323.170 ;
        RECT 2236.630 3143.590 2237.810 3144.770 ;
        RECT 2238.230 3143.590 2239.410 3144.770 ;
        RECT 2236.630 3141.990 2237.810 3143.170 ;
        RECT 2238.230 3141.990 2239.410 3143.170 ;
        RECT 2236.630 2963.590 2237.810 2964.770 ;
        RECT 2238.230 2963.590 2239.410 2964.770 ;
        RECT 2236.630 2961.990 2237.810 2963.170 ;
        RECT 2238.230 2961.990 2239.410 2963.170 ;
        RECT 2236.630 2783.590 2237.810 2784.770 ;
        RECT 2238.230 2783.590 2239.410 2784.770 ;
        RECT 2236.630 2781.990 2237.810 2783.170 ;
        RECT 2238.230 2781.990 2239.410 2783.170 ;
        RECT 2236.630 2603.590 2237.810 2604.770 ;
        RECT 2238.230 2603.590 2239.410 2604.770 ;
        RECT 2236.630 2601.990 2237.810 2603.170 ;
        RECT 2238.230 2601.990 2239.410 2603.170 ;
        RECT 2236.630 2423.590 2237.810 2424.770 ;
        RECT 2238.230 2423.590 2239.410 2424.770 ;
        RECT 2236.630 2421.990 2237.810 2423.170 ;
        RECT 2238.230 2421.990 2239.410 2423.170 ;
        RECT 2236.630 2243.590 2237.810 2244.770 ;
        RECT 2238.230 2243.590 2239.410 2244.770 ;
        RECT 2236.630 2241.990 2237.810 2243.170 ;
        RECT 2238.230 2241.990 2239.410 2243.170 ;
        RECT 2236.630 2063.590 2237.810 2064.770 ;
        RECT 2238.230 2063.590 2239.410 2064.770 ;
        RECT 2236.630 2061.990 2237.810 2063.170 ;
        RECT 2238.230 2061.990 2239.410 2063.170 ;
        RECT 2236.630 1883.590 2237.810 1884.770 ;
        RECT 2238.230 1883.590 2239.410 1884.770 ;
        RECT 2236.630 1881.990 2237.810 1883.170 ;
        RECT 2238.230 1881.990 2239.410 1883.170 ;
        RECT 2236.630 1703.590 2237.810 1704.770 ;
        RECT 2238.230 1703.590 2239.410 1704.770 ;
        RECT 2236.630 1701.990 2237.810 1703.170 ;
        RECT 2238.230 1701.990 2239.410 1703.170 ;
        RECT 2236.630 1523.590 2237.810 1524.770 ;
        RECT 2238.230 1523.590 2239.410 1524.770 ;
        RECT 2236.630 1521.990 2237.810 1523.170 ;
        RECT 2238.230 1521.990 2239.410 1523.170 ;
        RECT 2236.630 1343.590 2237.810 1344.770 ;
        RECT 2238.230 1343.590 2239.410 1344.770 ;
        RECT 2236.630 1341.990 2237.810 1343.170 ;
        RECT 2238.230 1341.990 2239.410 1343.170 ;
        RECT 2236.630 1163.590 2237.810 1164.770 ;
        RECT 2238.230 1163.590 2239.410 1164.770 ;
        RECT 2236.630 1161.990 2237.810 1163.170 ;
        RECT 2238.230 1161.990 2239.410 1163.170 ;
        RECT 2236.630 983.590 2237.810 984.770 ;
        RECT 2238.230 983.590 2239.410 984.770 ;
        RECT 2236.630 981.990 2237.810 983.170 ;
        RECT 2238.230 981.990 2239.410 983.170 ;
        RECT 2236.630 803.590 2237.810 804.770 ;
        RECT 2238.230 803.590 2239.410 804.770 ;
        RECT 2236.630 801.990 2237.810 803.170 ;
        RECT 2238.230 801.990 2239.410 803.170 ;
        RECT 2236.630 623.590 2237.810 624.770 ;
        RECT 2238.230 623.590 2239.410 624.770 ;
        RECT 2236.630 621.990 2237.810 623.170 ;
        RECT 2238.230 621.990 2239.410 623.170 ;
        RECT 2236.630 443.590 2237.810 444.770 ;
        RECT 2238.230 443.590 2239.410 444.770 ;
        RECT 2236.630 441.990 2237.810 443.170 ;
        RECT 2238.230 441.990 2239.410 443.170 ;
        RECT 2236.630 263.590 2237.810 264.770 ;
        RECT 2238.230 263.590 2239.410 264.770 ;
        RECT 2236.630 261.990 2237.810 263.170 ;
        RECT 2238.230 261.990 2239.410 263.170 ;
        RECT 2236.630 83.590 2237.810 84.770 ;
        RECT 2238.230 83.590 2239.410 84.770 ;
        RECT 2236.630 81.990 2237.810 83.170 ;
        RECT 2238.230 81.990 2239.410 83.170 ;
        RECT 2236.630 -18.860 2237.810 -17.680 ;
        RECT 2238.230 -18.860 2239.410 -17.680 ;
        RECT 2236.630 -20.460 2237.810 -19.280 ;
        RECT 2238.230 -20.460 2239.410 -19.280 ;
        RECT 2416.630 3538.960 2417.810 3540.140 ;
        RECT 2418.230 3538.960 2419.410 3540.140 ;
        RECT 2416.630 3537.360 2417.810 3538.540 ;
        RECT 2418.230 3537.360 2419.410 3538.540 ;
        RECT 2416.630 3503.590 2417.810 3504.770 ;
        RECT 2418.230 3503.590 2419.410 3504.770 ;
        RECT 2416.630 3501.990 2417.810 3503.170 ;
        RECT 2418.230 3501.990 2419.410 3503.170 ;
        RECT 2416.630 3323.590 2417.810 3324.770 ;
        RECT 2418.230 3323.590 2419.410 3324.770 ;
        RECT 2416.630 3321.990 2417.810 3323.170 ;
        RECT 2418.230 3321.990 2419.410 3323.170 ;
        RECT 2416.630 3143.590 2417.810 3144.770 ;
        RECT 2418.230 3143.590 2419.410 3144.770 ;
        RECT 2416.630 3141.990 2417.810 3143.170 ;
        RECT 2418.230 3141.990 2419.410 3143.170 ;
        RECT 2416.630 2963.590 2417.810 2964.770 ;
        RECT 2418.230 2963.590 2419.410 2964.770 ;
        RECT 2416.630 2961.990 2417.810 2963.170 ;
        RECT 2418.230 2961.990 2419.410 2963.170 ;
        RECT 2416.630 2783.590 2417.810 2784.770 ;
        RECT 2418.230 2783.590 2419.410 2784.770 ;
        RECT 2416.630 2781.990 2417.810 2783.170 ;
        RECT 2418.230 2781.990 2419.410 2783.170 ;
        RECT 2416.630 2603.590 2417.810 2604.770 ;
        RECT 2418.230 2603.590 2419.410 2604.770 ;
        RECT 2416.630 2601.990 2417.810 2603.170 ;
        RECT 2418.230 2601.990 2419.410 2603.170 ;
        RECT 2416.630 2423.590 2417.810 2424.770 ;
        RECT 2418.230 2423.590 2419.410 2424.770 ;
        RECT 2416.630 2421.990 2417.810 2423.170 ;
        RECT 2418.230 2421.990 2419.410 2423.170 ;
        RECT 2416.630 2243.590 2417.810 2244.770 ;
        RECT 2418.230 2243.590 2419.410 2244.770 ;
        RECT 2416.630 2241.990 2417.810 2243.170 ;
        RECT 2418.230 2241.990 2419.410 2243.170 ;
        RECT 2416.630 2063.590 2417.810 2064.770 ;
        RECT 2418.230 2063.590 2419.410 2064.770 ;
        RECT 2416.630 2061.990 2417.810 2063.170 ;
        RECT 2418.230 2061.990 2419.410 2063.170 ;
        RECT 2416.630 1883.590 2417.810 1884.770 ;
        RECT 2418.230 1883.590 2419.410 1884.770 ;
        RECT 2416.630 1881.990 2417.810 1883.170 ;
        RECT 2418.230 1881.990 2419.410 1883.170 ;
        RECT 2416.630 1703.590 2417.810 1704.770 ;
        RECT 2418.230 1703.590 2419.410 1704.770 ;
        RECT 2416.630 1701.990 2417.810 1703.170 ;
        RECT 2418.230 1701.990 2419.410 1703.170 ;
        RECT 2416.630 1523.590 2417.810 1524.770 ;
        RECT 2418.230 1523.590 2419.410 1524.770 ;
        RECT 2416.630 1521.990 2417.810 1523.170 ;
        RECT 2418.230 1521.990 2419.410 1523.170 ;
        RECT 2416.630 1343.590 2417.810 1344.770 ;
        RECT 2418.230 1343.590 2419.410 1344.770 ;
        RECT 2416.630 1341.990 2417.810 1343.170 ;
        RECT 2418.230 1341.990 2419.410 1343.170 ;
        RECT 2416.630 1163.590 2417.810 1164.770 ;
        RECT 2418.230 1163.590 2419.410 1164.770 ;
        RECT 2416.630 1161.990 2417.810 1163.170 ;
        RECT 2418.230 1161.990 2419.410 1163.170 ;
        RECT 2416.630 983.590 2417.810 984.770 ;
        RECT 2418.230 983.590 2419.410 984.770 ;
        RECT 2416.630 981.990 2417.810 983.170 ;
        RECT 2418.230 981.990 2419.410 983.170 ;
        RECT 2416.630 803.590 2417.810 804.770 ;
        RECT 2418.230 803.590 2419.410 804.770 ;
        RECT 2416.630 801.990 2417.810 803.170 ;
        RECT 2418.230 801.990 2419.410 803.170 ;
        RECT 2416.630 623.590 2417.810 624.770 ;
        RECT 2418.230 623.590 2419.410 624.770 ;
        RECT 2416.630 621.990 2417.810 623.170 ;
        RECT 2418.230 621.990 2419.410 623.170 ;
        RECT 2416.630 443.590 2417.810 444.770 ;
        RECT 2418.230 443.590 2419.410 444.770 ;
        RECT 2416.630 441.990 2417.810 443.170 ;
        RECT 2418.230 441.990 2419.410 443.170 ;
        RECT 2416.630 263.590 2417.810 264.770 ;
        RECT 2418.230 263.590 2419.410 264.770 ;
        RECT 2416.630 261.990 2417.810 263.170 ;
        RECT 2418.230 261.990 2419.410 263.170 ;
        RECT 2416.630 83.590 2417.810 84.770 ;
        RECT 2418.230 83.590 2419.410 84.770 ;
        RECT 2416.630 81.990 2417.810 83.170 ;
        RECT 2418.230 81.990 2419.410 83.170 ;
        RECT 2416.630 -18.860 2417.810 -17.680 ;
        RECT 2418.230 -18.860 2419.410 -17.680 ;
        RECT 2416.630 -20.460 2417.810 -19.280 ;
        RECT 2418.230 -20.460 2419.410 -19.280 ;
        RECT 2596.630 3538.960 2597.810 3540.140 ;
        RECT 2598.230 3538.960 2599.410 3540.140 ;
        RECT 2596.630 3537.360 2597.810 3538.540 ;
        RECT 2598.230 3537.360 2599.410 3538.540 ;
        RECT 2596.630 3503.590 2597.810 3504.770 ;
        RECT 2598.230 3503.590 2599.410 3504.770 ;
        RECT 2596.630 3501.990 2597.810 3503.170 ;
        RECT 2598.230 3501.990 2599.410 3503.170 ;
        RECT 2596.630 3323.590 2597.810 3324.770 ;
        RECT 2598.230 3323.590 2599.410 3324.770 ;
        RECT 2596.630 3321.990 2597.810 3323.170 ;
        RECT 2598.230 3321.990 2599.410 3323.170 ;
        RECT 2596.630 3143.590 2597.810 3144.770 ;
        RECT 2598.230 3143.590 2599.410 3144.770 ;
        RECT 2596.630 3141.990 2597.810 3143.170 ;
        RECT 2598.230 3141.990 2599.410 3143.170 ;
        RECT 2596.630 2963.590 2597.810 2964.770 ;
        RECT 2598.230 2963.590 2599.410 2964.770 ;
        RECT 2596.630 2961.990 2597.810 2963.170 ;
        RECT 2598.230 2961.990 2599.410 2963.170 ;
        RECT 2596.630 2783.590 2597.810 2784.770 ;
        RECT 2598.230 2783.590 2599.410 2784.770 ;
        RECT 2596.630 2781.990 2597.810 2783.170 ;
        RECT 2598.230 2781.990 2599.410 2783.170 ;
        RECT 2596.630 2603.590 2597.810 2604.770 ;
        RECT 2598.230 2603.590 2599.410 2604.770 ;
        RECT 2596.630 2601.990 2597.810 2603.170 ;
        RECT 2598.230 2601.990 2599.410 2603.170 ;
        RECT 2596.630 2423.590 2597.810 2424.770 ;
        RECT 2598.230 2423.590 2599.410 2424.770 ;
        RECT 2596.630 2421.990 2597.810 2423.170 ;
        RECT 2598.230 2421.990 2599.410 2423.170 ;
        RECT 2596.630 2243.590 2597.810 2244.770 ;
        RECT 2598.230 2243.590 2599.410 2244.770 ;
        RECT 2596.630 2241.990 2597.810 2243.170 ;
        RECT 2598.230 2241.990 2599.410 2243.170 ;
        RECT 2596.630 2063.590 2597.810 2064.770 ;
        RECT 2598.230 2063.590 2599.410 2064.770 ;
        RECT 2596.630 2061.990 2597.810 2063.170 ;
        RECT 2598.230 2061.990 2599.410 2063.170 ;
        RECT 2596.630 1883.590 2597.810 1884.770 ;
        RECT 2598.230 1883.590 2599.410 1884.770 ;
        RECT 2596.630 1881.990 2597.810 1883.170 ;
        RECT 2598.230 1881.990 2599.410 1883.170 ;
        RECT 2596.630 1703.590 2597.810 1704.770 ;
        RECT 2598.230 1703.590 2599.410 1704.770 ;
        RECT 2596.630 1701.990 2597.810 1703.170 ;
        RECT 2598.230 1701.990 2599.410 1703.170 ;
        RECT 2596.630 1523.590 2597.810 1524.770 ;
        RECT 2598.230 1523.590 2599.410 1524.770 ;
        RECT 2596.630 1521.990 2597.810 1523.170 ;
        RECT 2598.230 1521.990 2599.410 1523.170 ;
        RECT 2596.630 1343.590 2597.810 1344.770 ;
        RECT 2598.230 1343.590 2599.410 1344.770 ;
        RECT 2596.630 1341.990 2597.810 1343.170 ;
        RECT 2598.230 1341.990 2599.410 1343.170 ;
        RECT 2596.630 1163.590 2597.810 1164.770 ;
        RECT 2598.230 1163.590 2599.410 1164.770 ;
        RECT 2596.630 1161.990 2597.810 1163.170 ;
        RECT 2598.230 1161.990 2599.410 1163.170 ;
        RECT 2596.630 983.590 2597.810 984.770 ;
        RECT 2598.230 983.590 2599.410 984.770 ;
        RECT 2596.630 981.990 2597.810 983.170 ;
        RECT 2598.230 981.990 2599.410 983.170 ;
        RECT 2596.630 803.590 2597.810 804.770 ;
        RECT 2598.230 803.590 2599.410 804.770 ;
        RECT 2596.630 801.990 2597.810 803.170 ;
        RECT 2598.230 801.990 2599.410 803.170 ;
        RECT 2596.630 623.590 2597.810 624.770 ;
        RECT 2598.230 623.590 2599.410 624.770 ;
        RECT 2596.630 621.990 2597.810 623.170 ;
        RECT 2598.230 621.990 2599.410 623.170 ;
        RECT 2596.630 443.590 2597.810 444.770 ;
        RECT 2598.230 443.590 2599.410 444.770 ;
        RECT 2596.630 441.990 2597.810 443.170 ;
        RECT 2598.230 441.990 2599.410 443.170 ;
        RECT 2596.630 263.590 2597.810 264.770 ;
        RECT 2598.230 263.590 2599.410 264.770 ;
        RECT 2596.630 261.990 2597.810 263.170 ;
        RECT 2598.230 261.990 2599.410 263.170 ;
        RECT 2596.630 83.590 2597.810 84.770 ;
        RECT 2598.230 83.590 2599.410 84.770 ;
        RECT 2596.630 81.990 2597.810 83.170 ;
        RECT 2598.230 81.990 2599.410 83.170 ;
        RECT 2596.630 -18.860 2597.810 -17.680 ;
        RECT 2598.230 -18.860 2599.410 -17.680 ;
        RECT 2596.630 -20.460 2597.810 -19.280 ;
        RECT 2598.230 -20.460 2599.410 -19.280 ;
        RECT 2776.630 3538.960 2777.810 3540.140 ;
        RECT 2778.230 3538.960 2779.410 3540.140 ;
        RECT 2776.630 3537.360 2777.810 3538.540 ;
        RECT 2778.230 3537.360 2779.410 3538.540 ;
        RECT 2776.630 3503.590 2777.810 3504.770 ;
        RECT 2778.230 3503.590 2779.410 3504.770 ;
        RECT 2776.630 3501.990 2777.810 3503.170 ;
        RECT 2778.230 3501.990 2779.410 3503.170 ;
        RECT 2776.630 3323.590 2777.810 3324.770 ;
        RECT 2778.230 3323.590 2779.410 3324.770 ;
        RECT 2776.630 3321.990 2777.810 3323.170 ;
        RECT 2778.230 3321.990 2779.410 3323.170 ;
        RECT 2776.630 3143.590 2777.810 3144.770 ;
        RECT 2778.230 3143.590 2779.410 3144.770 ;
        RECT 2776.630 3141.990 2777.810 3143.170 ;
        RECT 2778.230 3141.990 2779.410 3143.170 ;
        RECT 2776.630 2963.590 2777.810 2964.770 ;
        RECT 2778.230 2963.590 2779.410 2964.770 ;
        RECT 2776.630 2961.990 2777.810 2963.170 ;
        RECT 2778.230 2961.990 2779.410 2963.170 ;
        RECT 2776.630 2783.590 2777.810 2784.770 ;
        RECT 2778.230 2783.590 2779.410 2784.770 ;
        RECT 2776.630 2781.990 2777.810 2783.170 ;
        RECT 2778.230 2781.990 2779.410 2783.170 ;
        RECT 2776.630 2603.590 2777.810 2604.770 ;
        RECT 2778.230 2603.590 2779.410 2604.770 ;
        RECT 2776.630 2601.990 2777.810 2603.170 ;
        RECT 2778.230 2601.990 2779.410 2603.170 ;
        RECT 2776.630 2423.590 2777.810 2424.770 ;
        RECT 2778.230 2423.590 2779.410 2424.770 ;
        RECT 2776.630 2421.990 2777.810 2423.170 ;
        RECT 2778.230 2421.990 2779.410 2423.170 ;
        RECT 2776.630 2243.590 2777.810 2244.770 ;
        RECT 2778.230 2243.590 2779.410 2244.770 ;
        RECT 2776.630 2241.990 2777.810 2243.170 ;
        RECT 2778.230 2241.990 2779.410 2243.170 ;
        RECT 2776.630 2063.590 2777.810 2064.770 ;
        RECT 2778.230 2063.590 2779.410 2064.770 ;
        RECT 2776.630 2061.990 2777.810 2063.170 ;
        RECT 2778.230 2061.990 2779.410 2063.170 ;
        RECT 2776.630 1883.590 2777.810 1884.770 ;
        RECT 2778.230 1883.590 2779.410 1884.770 ;
        RECT 2776.630 1881.990 2777.810 1883.170 ;
        RECT 2778.230 1881.990 2779.410 1883.170 ;
        RECT 2776.630 1703.590 2777.810 1704.770 ;
        RECT 2778.230 1703.590 2779.410 1704.770 ;
        RECT 2776.630 1701.990 2777.810 1703.170 ;
        RECT 2778.230 1701.990 2779.410 1703.170 ;
        RECT 2776.630 1523.590 2777.810 1524.770 ;
        RECT 2778.230 1523.590 2779.410 1524.770 ;
        RECT 2776.630 1521.990 2777.810 1523.170 ;
        RECT 2778.230 1521.990 2779.410 1523.170 ;
        RECT 2776.630 1343.590 2777.810 1344.770 ;
        RECT 2778.230 1343.590 2779.410 1344.770 ;
        RECT 2776.630 1341.990 2777.810 1343.170 ;
        RECT 2778.230 1341.990 2779.410 1343.170 ;
        RECT 2776.630 1163.590 2777.810 1164.770 ;
        RECT 2778.230 1163.590 2779.410 1164.770 ;
        RECT 2776.630 1161.990 2777.810 1163.170 ;
        RECT 2778.230 1161.990 2779.410 1163.170 ;
        RECT 2776.630 983.590 2777.810 984.770 ;
        RECT 2778.230 983.590 2779.410 984.770 ;
        RECT 2776.630 981.990 2777.810 983.170 ;
        RECT 2778.230 981.990 2779.410 983.170 ;
        RECT 2776.630 803.590 2777.810 804.770 ;
        RECT 2778.230 803.590 2779.410 804.770 ;
        RECT 2776.630 801.990 2777.810 803.170 ;
        RECT 2778.230 801.990 2779.410 803.170 ;
        RECT 2776.630 623.590 2777.810 624.770 ;
        RECT 2778.230 623.590 2779.410 624.770 ;
        RECT 2776.630 621.990 2777.810 623.170 ;
        RECT 2778.230 621.990 2779.410 623.170 ;
        RECT 2776.630 443.590 2777.810 444.770 ;
        RECT 2778.230 443.590 2779.410 444.770 ;
        RECT 2776.630 441.990 2777.810 443.170 ;
        RECT 2778.230 441.990 2779.410 443.170 ;
        RECT 2776.630 263.590 2777.810 264.770 ;
        RECT 2778.230 263.590 2779.410 264.770 ;
        RECT 2776.630 261.990 2777.810 263.170 ;
        RECT 2778.230 261.990 2779.410 263.170 ;
        RECT 2776.630 83.590 2777.810 84.770 ;
        RECT 2778.230 83.590 2779.410 84.770 ;
        RECT 2776.630 81.990 2777.810 83.170 ;
        RECT 2778.230 81.990 2779.410 83.170 ;
        RECT 2776.630 -18.860 2777.810 -17.680 ;
        RECT 2778.230 -18.860 2779.410 -17.680 ;
        RECT 2776.630 -20.460 2777.810 -19.280 ;
        RECT 2778.230 -20.460 2779.410 -19.280 ;
        RECT 2942.660 3538.960 2943.840 3540.140 ;
        RECT 2944.260 3538.960 2945.440 3540.140 ;
        RECT 2942.660 3537.360 2943.840 3538.540 ;
        RECT 2944.260 3537.360 2945.440 3538.540 ;
        RECT 2942.660 3503.590 2943.840 3504.770 ;
        RECT 2944.260 3503.590 2945.440 3504.770 ;
        RECT 2942.660 3501.990 2943.840 3503.170 ;
        RECT 2944.260 3501.990 2945.440 3503.170 ;
        RECT 2942.660 3323.590 2943.840 3324.770 ;
        RECT 2944.260 3323.590 2945.440 3324.770 ;
        RECT 2942.660 3321.990 2943.840 3323.170 ;
        RECT 2944.260 3321.990 2945.440 3323.170 ;
        RECT 2942.660 3143.590 2943.840 3144.770 ;
        RECT 2944.260 3143.590 2945.440 3144.770 ;
        RECT 2942.660 3141.990 2943.840 3143.170 ;
        RECT 2944.260 3141.990 2945.440 3143.170 ;
        RECT 2942.660 2963.590 2943.840 2964.770 ;
        RECT 2944.260 2963.590 2945.440 2964.770 ;
        RECT 2942.660 2961.990 2943.840 2963.170 ;
        RECT 2944.260 2961.990 2945.440 2963.170 ;
        RECT 2942.660 2783.590 2943.840 2784.770 ;
        RECT 2944.260 2783.590 2945.440 2784.770 ;
        RECT 2942.660 2781.990 2943.840 2783.170 ;
        RECT 2944.260 2781.990 2945.440 2783.170 ;
        RECT 2942.660 2603.590 2943.840 2604.770 ;
        RECT 2944.260 2603.590 2945.440 2604.770 ;
        RECT 2942.660 2601.990 2943.840 2603.170 ;
        RECT 2944.260 2601.990 2945.440 2603.170 ;
        RECT 2942.660 2423.590 2943.840 2424.770 ;
        RECT 2944.260 2423.590 2945.440 2424.770 ;
        RECT 2942.660 2421.990 2943.840 2423.170 ;
        RECT 2944.260 2421.990 2945.440 2423.170 ;
        RECT 2942.660 2243.590 2943.840 2244.770 ;
        RECT 2944.260 2243.590 2945.440 2244.770 ;
        RECT 2942.660 2241.990 2943.840 2243.170 ;
        RECT 2944.260 2241.990 2945.440 2243.170 ;
        RECT 2942.660 2063.590 2943.840 2064.770 ;
        RECT 2944.260 2063.590 2945.440 2064.770 ;
        RECT 2942.660 2061.990 2943.840 2063.170 ;
        RECT 2944.260 2061.990 2945.440 2063.170 ;
        RECT 2942.660 1883.590 2943.840 1884.770 ;
        RECT 2944.260 1883.590 2945.440 1884.770 ;
        RECT 2942.660 1881.990 2943.840 1883.170 ;
        RECT 2944.260 1881.990 2945.440 1883.170 ;
        RECT 2942.660 1703.590 2943.840 1704.770 ;
        RECT 2944.260 1703.590 2945.440 1704.770 ;
        RECT 2942.660 1701.990 2943.840 1703.170 ;
        RECT 2944.260 1701.990 2945.440 1703.170 ;
        RECT 2942.660 1523.590 2943.840 1524.770 ;
        RECT 2944.260 1523.590 2945.440 1524.770 ;
        RECT 2942.660 1521.990 2943.840 1523.170 ;
        RECT 2944.260 1521.990 2945.440 1523.170 ;
        RECT 2942.660 1343.590 2943.840 1344.770 ;
        RECT 2944.260 1343.590 2945.440 1344.770 ;
        RECT 2942.660 1341.990 2943.840 1343.170 ;
        RECT 2944.260 1341.990 2945.440 1343.170 ;
        RECT 2942.660 1163.590 2943.840 1164.770 ;
        RECT 2944.260 1163.590 2945.440 1164.770 ;
        RECT 2942.660 1161.990 2943.840 1163.170 ;
        RECT 2944.260 1161.990 2945.440 1163.170 ;
        RECT 2942.660 983.590 2943.840 984.770 ;
        RECT 2944.260 983.590 2945.440 984.770 ;
        RECT 2942.660 981.990 2943.840 983.170 ;
        RECT 2944.260 981.990 2945.440 983.170 ;
        RECT 2942.660 803.590 2943.840 804.770 ;
        RECT 2944.260 803.590 2945.440 804.770 ;
        RECT 2942.660 801.990 2943.840 803.170 ;
        RECT 2944.260 801.990 2945.440 803.170 ;
        RECT 2942.660 623.590 2943.840 624.770 ;
        RECT 2944.260 623.590 2945.440 624.770 ;
        RECT 2942.660 621.990 2943.840 623.170 ;
        RECT 2944.260 621.990 2945.440 623.170 ;
        RECT 2942.660 443.590 2943.840 444.770 ;
        RECT 2944.260 443.590 2945.440 444.770 ;
        RECT 2942.660 441.990 2943.840 443.170 ;
        RECT 2944.260 441.990 2945.440 443.170 ;
        RECT 2942.660 263.590 2943.840 264.770 ;
        RECT 2944.260 263.590 2945.440 264.770 ;
        RECT 2942.660 261.990 2943.840 263.170 ;
        RECT 2944.260 261.990 2945.440 263.170 ;
        RECT 2942.660 83.590 2943.840 84.770 ;
        RECT 2944.260 83.590 2945.440 84.770 ;
        RECT 2942.660 81.990 2943.840 83.170 ;
        RECT 2944.260 81.990 2945.440 83.170 ;
        RECT 2942.660 -18.860 2943.840 -17.680 ;
        RECT 2944.260 -18.860 2945.440 -17.680 ;
        RECT 2942.660 -20.460 2943.840 -19.280 ;
        RECT 2944.260 -20.460 2945.440 -19.280 ;
      LAYER met5 ;
        RECT -25.980 3537.200 2945.600 3540.300 ;
        RECT -45.180 3501.830 2964.800 3504.930 ;
        RECT -45.180 3321.830 2964.800 3324.930 ;
        RECT -45.180 3141.830 2964.800 3144.930 ;
        RECT -45.180 2961.830 2964.800 2964.930 ;
        RECT -45.180 2781.830 2964.800 2784.930 ;
        RECT -45.180 2601.830 2964.800 2604.930 ;
        RECT -45.180 2421.830 2964.800 2424.930 ;
        RECT -45.180 2241.830 2964.800 2244.930 ;
        RECT -45.180 2061.830 2964.800 2064.930 ;
        RECT -45.180 1881.830 2964.800 1884.930 ;
        RECT -45.180 1701.830 2964.800 1704.930 ;
        RECT -45.180 1521.830 2964.800 1524.930 ;
        RECT -45.180 1341.830 2964.800 1344.930 ;
        RECT -45.180 1161.830 2964.800 1164.930 ;
        RECT -45.180 981.830 2964.800 984.930 ;
        RECT -45.180 801.830 2964.800 804.930 ;
        RECT -45.180 621.830 2964.800 624.930 ;
        RECT -45.180 441.830 2964.800 444.930 ;
        RECT -45.180 261.830 2964.800 264.930 ;
        RECT -45.180 81.830 2964.800 84.930 ;
        RECT -25.980 -20.620 2945.600 -17.520 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 -4.800 110.450 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.630 473.520 407.950 473.580 ;
        RECT 412.230 473.520 412.550 473.580 ;
        RECT 407.630 473.380 412.550 473.520 ;
        RECT 407.630 473.320 407.950 473.380 ;
        RECT 412.230 473.320 412.550 473.380 ;
        RECT 115.530 24.040 115.850 24.100 ;
        RECT 407.630 24.040 407.950 24.100 ;
        RECT 115.530 23.900 407.950 24.040 ;
        RECT 115.530 23.840 115.850 23.900 ;
        RECT 407.630 23.840 407.950 23.900 ;
      LAYER via ;
        RECT 407.660 473.320 407.920 473.580 ;
        RECT 412.260 473.320 412.520 473.580 ;
        RECT 115.560 23.840 115.820 24.100 ;
        RECT 407.660 23.840 407.920 24.100 ;
      LAYER met2 ;
        RECT 412.510 500.000 412.790 504.000 ;
        RECT 412.550 498.850 412.690 500.000 ;
        RECT 412.320 498.710 412.690 498.850 ;
        RECT 412.320 473.610 412.460 498.710 ;
        RECT 407.660 473.290 407.920 473.610 ;
        RECT 412.260 473.290 412.520 473.610 ;
        RECT 407.720 24.130 407.860 473.290 ;
        RECT 115.560 23.810 115.820 24.130 ;
        RECT 407.660 23.810 407.920 24.130 ;
        RECT 115.620 2.400 115.760 23.810 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.090 499.360 408.410 499.420 ;
        RECT 412.920 499.360 413.240 499.420 ;
        RECT 408.090 499.220 413.240 499.360 ;
        RECT 408.090 499.160 408.410 499.220 ;
        RECT 412.920 499.160 413.240 499.220 ;
        RECT 121.050 24.380 121.370 24.440 ;
        RECT 408.090 24.380 408.410 24.440 ;
        RECT 121.050 24.240 408.410 24.380 ;
        RECT 121.050 24.180 121.370 24.240 ;
        RECT 408.090 24.180 408.410 24.240 ;
      LAYER via ;
        RECT 408.120 499.160 408.380 499.420 ;
        RECT 412.950 499.160 413.210 499.420 ;
        RECT 121.080 24.180 121.340 24.440 ;
        RECT 408.120 24.180 408.380 24.440 ;
      LAYER met2 ;
        RECT 412.970 500.000 413.250 504.000 ;
        RECT 413.010 499.450 413.150 500.000 ;
        RECT 408.120 499.130 408.380 499.450 ;
        RECT 412.950 499.130 413.210 499.450 ;
        RECT 408.180 24.470 408.320 499.130 ;
        RECT 121.080 24.150 121.340 24.470 ;
        RECT 408.120 24.150 408.380 24.470 ;
        RECT 121.140 2.400 121.280 24.150 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.990 17.240 415.310 17.300 ;
        RECT 179.330 17.100 415.310 17.240 ;
        RECT 143.130 16.900 143.450 16.960 ;
        RECT 179.330 16.900 179.470 17.100 ;
        RECT 414.990 17.040 415.310 17.100 ;
        RECT 143.130 16.760 179.470 16.900 ;
        RECT 143.130 16.700 143.450 16.760 ;
      LAYER via ;
        RECT 143.160 16.700 143.420 16.960 ;
        RECT 415.020 17.040 415.280 17.300 ;
      LAYER met2 ;
        RECT 414.810 500.000 415.090 504.000 ;
        RECT 414.850 498.850 414.990 500.000 ;
        RECT 414.850 498.710 415.220 498.850 ;
        RECT 415.080 17.330 415.220 498.710 ;
        RECT 415.020 17.010 415.280 17.330 ;
        RECT 143.160 16.670 143.420 16.990 ;
        RECT 143.220 2.400 143.360 16.670 ;
        RECT 143.010 -4.800 143.570 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.790 487.460 429.110 487.520 ;
        RECT 430.630 487.460 430.950 487.520 ;
        RECT 428.790 487.320 430.950 487.460 ;
        RECT 428.790 487.260 429.110 487.320 ;
        RECT 430.630 487.260 430.950 487.320 ;
        RECT 330.810 18.940 331.130 19.000 ;
        RECT 428.790 18.940 429.110 19.000 ;
        RECT 330.810 18.800 429.110 18.940 ;
        RECT 330.810 18.740 331.130 18.800 ;
        RECT 428.790 18.740 429.110 18.800 ;
      LAYER via ;
        RECT 428.820 487.260 429.080 487.520 ;
        RECT 430.660 487.260 430.920 487.520 ;
        RECT 330.840 18.740 331.100 19.000 ;
        RECT 428.820 18.740 429.080 19.000 ;
      LAYER met2 ;
        RECT 430.450 500.000 430.730 504.000 ;
        RECT 430.490 499.020 430.630 500.000 ;
        RECT 430.490 498.880 430.860 499.020 ;
        RECT 430.720 487.550 430.860 498.880 ;
        RECT 428.820 487.230 429.080 487.550 ;
        RECT 430.660 487.230 430.920 487.550 ;
        RECT 428.880 19.030 429.020 487.230 ;
        RECT 330.840 18.710 331.100 19.030 ;
        RECT 428.820 18.710 429.080 19.030 ;
        RECT 330.900 2.400 331.040 18.710 ;
        RECT 330.690 -4.800 331.250 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 347.370 19.280 347.690 19.340 ;
        RECT 432.930 19.280 433.250 19.340 ;
        RECT 347.370 19.140 433.250 19.280 ;
        RECT 347.370 19.080 347.690 19.140 ;
        RECT 432.930 19.080 433.250 19.140 ;
      LAYER via ;
        RECT 347.400 19.080 347.660 19.340 ;
        RECT 432.960 19.080 433.220 19.340 ;
      LAYER met2 ;
        RECT 431.830 500.000 432.110 504.000 ;
        RECT 431.870 499.645 432.010 500.000 ;
        RECT 431.800 499.275 432.080 499.645 ;
        RECT 432.490 491.115 432.770 491.485 ;
        RECT 432.560 448.570 432.700 491.115 ;
        RECT 432.560 448.430 433.160 448.570 ;
        RECT 433.020 19.370 433.160 448.430 ;
        RECT 347.400 19.050 347.660 19.370 ;
        RECT 432.960 19.050 433.220 19.370 ;
        RECT 347.460 2.400 347.600 19.050 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 431.800 499.320 432.080 499.600 ;
        RECT 432.490 491.160 432.770 491.440 ;
      LAYER met3 ;
        RECT 431.775 499.620 432.105 499.625 ;
        RECT 431.750 499.610 432.130 499.620 ;
        RECT 431.320 499.310 432.130 499.610 ;
        RECT 431.750 499.300 432.130 499.310 ;
        RECT 431.775 499.295 432.105 499.300 ;
        RECT 431.750 491.450 432.130 491.460 ;
        RECT 432.465 491.450 432.795 491.465 ;
        RECT 431.750 491.150 432.795 491.450 ;
        RECT 431.750 491.140 432.130 491.150 ;
        RECT 432.465 491.135 432.795 491.150 ;
      LAYER via3 ;
        RECT 431.780 499.300 432.100 499.620 ;
        RECT 431.780 491.140 432.100 491.460 ;
      LAYER met4 ;
        RECT 431.775 499.295 432.105 499.625 ;
        RECT 431.790 491.465 432.090 499.295 ;
        RECT 431.775 491.135 432.105 491.465 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 433.160 500.520 433.480 500.780 ;
        RECT 433.250 500.040 433.390 500.520 ;
        RECT 433.250 499.900 434.540 500.040 ;
        RECT 433.390 497.320 433.710 497.380 ;
        RECT 434.400 497.320 434.540 499.900 ;
        RECT 433.390 497.180 434.540 497.320 ;
        RECT 433.390 497.120 433.710 497.180 ;
        RECT 363.930 19.620 364.250 19.680 ;
        RECT 433.390 19.620 433.710 19.680 ;
        RECT 363.930 19.480 433.710 19.620 ;
        RECT 363.930 19.420 364.250 19.480 ;
        RECT 433.390 19.420 433.710 19.480 ;
      LAYER via ;
        RECT 433.190 500.520 433.450 500.780 ;
        RECT 433.420 497.120 433.680 497.380 ;
        RECT 363.960 19.420 364.220 19.680 ;
        RECT 433.420 19.420 433.680 19.680 ;
      LAYER met2 ;
        RECT 433.210 500.810 433.490 504.000 ;
        RECT 433.190 500.490 433.490 500.810 ;
        RECT 433.210 500.000 433.490 500.490 ;
        RECT 433.420 497.090 433.680 497.410 ;
        RECT 433.480 19.710 433.620 497.090 ;
        RECT 363.960 19.390 364.220 19.710 ;
        RECT 433.420 19.390 433.680 19.710 ;
        RECT 364.020 2.400 364.160 19.390 ;
        RECT 363.810 -4.800 364.370 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 472.840 435.090 472.900 ;
        RECT 437.990 472.840 438.310 472.900 ;
        RECT 434.770 472.700 438.310 472.840 ;
        RECT 434.770 472.640 435.090 472.700 ;
        RECT 437.990 472.640 438.310 472.700 ;
        RECT 380.490 19.960 380.810 20.020 ;
        RECT 437.990 19.960 438.310 20.020 ;
        RECT 380.490 19.820 438.310 19.960 ;
        RECT 380.490 19.760 380.810 19.820 ;
        RECT 437.990 19.760 438.310 19.820 ;
      LAYER via ;
        RECT 434.800 472.640 435.060 472.900 ;
        RECT 438.020 472.640 438.280 472.900 ;
        RECT 380.520 19.760 380.780 20.020 ;
        RECT 438.020 19.760 438.280 20.020 ;
      LAYER met2 ;
        RECT 434.590 500.000 434.870 504.000 ;
        RECT 434.630 498.680 434.770 500.000 ;
        RECT 434.630 498.540 435.000 498.680 ;
        RECT 434.860 472.930 435.000 498.540 ;
        RECT 434.800 472.610 435.060 472.930 ;
        RECT 438.020 472.610 438.280 472.930 ;
        RECT 438.080 20.050 438.220 472.610 ;
        RECT 380.520 19.730 380.780 20.050 ;
        RECT 438.020 19.730 438.280 20.050 ;
        RECT 380.580 2.400 380.720 19.730 ;
        RECT 380.370 -4.800 380.930 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.920 498.820 436.240 499.080 ;
        RECT 436.010 498.060 436.150 498.820 ;
        RECT 435.690 497.860 436.150 498.060 ;
        RECT 435.690 497.800 436.010 497.860 ;
        RECT 436.150 473.520 436.470 473.580 ;
        RECT 437.530 473.520 437.850 473.580 ;
        RECT 436.150 473.380 437.850 473.520 ;
        RECT 436.150 473.320 436.470 473.380 ;
        RECT 437.530 473.320 437.850 473.380 ;
        RECT 397.050 20.300 397.370 20.360 ;
        RECT 437.530 20.300 437.850 20.360 ;
        RECT 397.050 20.160 437.850 20.300 ;
        RECT 397.050 20.100 397.370 20.160 ;
        RECT 437.530 20.100 437.850 20.160 ;
      LAYER via ;
        RECT 435.950 498.820 436.210 499.080 ;
        RECT 435.720 497.800 435.980 498.060 ;
        RECT 436.180 473.320 436.440 473.580 ;
        RECT 437.560 473.320 437.820 473.580 ;
        RECT 397.080 20.100 397.340 20.360 ;
        RECT 437.560 20.100 437.820 20.360 ;
      LAYER met2 ;
        RECT 435.970 500.000 436.250 504.000 ;
        RECT 436.010 499.110 436.150 500.000 ;
        RECT 435.950 498.790 436.210 499.110 ;
        RECT 435.720 498.000 435.980 498.090 ;
        RECT 435.720 497.860 436.380 498.000 ;
        RECT 435.720 497.770 435.980 497.860 ;
        RECT 436.240 473.610 436.380 497.860 ;
        RECT 436.180 473.290 436.440 473.610 ;
        RECT 437.560 473.290 437.820 473.610 ;
        RECT 437.620 20.390 437.760 473.290 ;
        RECT 397.080 20.070 397.340 20.390 ;
        RECT 437.560 20.070 437.820 20.390 ;
        RECT 397.140 2.400 397.280 20.070 ;
        RECT 396.930 -4.800 397.490 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.610 17.920 436.930 17.980 ;
        RECT 420.830 17.780 436.930 17.920 ;
        RECT 413.610 17.580 413.930 17.640 ;
        RECT 420.830 17.580 420.970 17.780 ;
        RECT 436.610 17.720 436.930 17.780 ;
        RECT 413.610 17.440 420.970 17.580 ;
        RECT 413.610 17.380 413.930 17.440 ;
      LAYER via ;
        RECT 413.640 17.380 413.900 17.640 ;
        RECT 436.640 17.720 436.900 17.980 ;
      LAYER met2 ;
        RECT 437.350 500.000 437.630 504.000 ;
        RECT 437.390 499.645 437.530 500.000 ;
        RECT 437.320 499.275 437.600 499.645 ;
        RECT 436.630 497.235 436.910 497.605 ;
        RECT 436.700 18.010 436.840 497.235 ;
        RECT 436.640 17.690 436.900 18.010 ;
        RECT 413.640 17.350 413.900 17.670 ;
        RECT 413.700 2.400 413.840 17.350 ;
        RECT 413.490 -4.800 414.050 2.400 ;
      LAYER via2 ;
        RECT 437.320 499.320 437.600 499.600 ;
        RECT 436.630 497.280 436.910 497.560 ;
      LAYER met3 ;
        RECT 437.295 499.610 437.625 499.625 ;
        RECT 436.390 499.310 437.625 499.610 ;
        RECT 436.390 497.585 436.690 499.310 ;
        RECT 437.295 499.295 437.625 499.310 ;
        RECT 436.390 497.270 436.935 497.585 ;
        RECT 436.605 497.255 436.935 497.270 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 438.910 497.800 439.230 498.060 ;
        RECT 435.230 496.640 435.550 496.700 ;
        RECT 439.000 496.640 439.140 497.800 ;
        RECT 435.230 496.500 439.140 496.640 ;
        RECT 435.230 496.440 435.550 496.500 ;
        RECT 430.170 17.580 430.490 17.640 ;
        RECT 436.150 17.580 436.470 17.640 ;
        RECT 430.170 17.440 436.470 17.580 ;
        RECT 430.170 17.380 430.490 17.440 ;
        RECT 436.150 17.380 436.470 17.440 ;
      LAYER via ;
        RECT 438.940 497.800 439.200 498.060 ;
        RECT 435.260 496.440 435.520 496.700 ;
        RECT 430.200 17.380 430.460 17.640 ;
        RECT 436.180 17.380 436.440 17.640 ;
      LAYER met2 ;
        RECT 438.730 500.000 439.010 504.000 ;
        RECT 438.770 498.850 438.910 500.000 ;
        RECT 438.770 498.710 439.140 498.850 ;
        RECT 439.000 498.090 439.140 498.710 ;
        RECT 438.940 497.770 439.200 498.090 ;
        RECT 435.260 496.410 435.520 496.730 ;
        RECT 435.320 472.840 435.460 496.410 ;
        RECT 435.320 472.700 436.380 472.840 ;
        RECT 436.240 17.670 436.380 472.700 ;
        RECT 430.200 17.350 430.460 17.670 ;
        RECT 436.180 17.350 436.440 17.670 ;
        RECT 430.260 2.400 430.400 17.350 ;
        RECT 430.050 -4.800 430.610 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 440.060 499.500 440.380 499.760 ;
        RECT 439.370 497.660 439.690 497.720 ;
        RECT 440.150 497.660 440.290 499.500 ;
        RECT 439.370 497.520 440.290 497.660 ;
        RECT 439.370 497.460 439.690 497.520 ;
        RECT 435.690 472.160 436.010 472.220 ;
        RECT 439.370 472.160 439.690 472.220 ;
        RECT 435.690 472.020 439.690 472.160 ;
        RECT 435.690 471.960 436.010 472.020 ;
        RECT 439.370 471.960 439.690 472.020 ;
        RECT 435.690 15.880 436.010 15.940 ;
        RECT 446.730 15.880 447.050 15.940 ;
        RECT 435.690 15.740 447.050 15.880 ;
        RECT 435.690 15.680 436.010 15.740 ;
        RECT 446.730 15.680 447.050 15.740 ;
      LAYER via ;
        RECT 440.090 499.500 440.350 499.760 ;
        RECT 439.400 497.460 439.660 497.720 ;
        RECT 435.720 471.960 435.980 472.220 ;
        RECT 439.400 471.960 439.660 472.220 ;
        RECT 435.720 15.680 435.980 15.940 ;
        RECT 446.760 15.680 447.020 15.940 ;
      LAYER met2 ;
        RECT 440.110 500.000 440.390 504.000 ;
        RECT 440.150 499.790 440.290 500.000 ;
        RECT 440.090 499.470 440.350 499.790 ;
        RECT 439.400 497.430 439.660 497.750 ;
        RECT 439.460 472.250 439.600 497.430 ;
        RECT 435.720 471.930 435.980 472.250 ;
        RECT 439.400 471.930 439.660 472.250 ;
        RECT 435.780 15.970 435.920 471.930 ;
        RECT 435.720 15.650 435.980 15.970 ;
        RECT 446.760 15.650 447.020 15.970 ;
        RECT 446.820 2.400 446.960 15.650 ;
        RECT 446.610 -4.800 447.170 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.440 499.160 441.760 499.420 ;
        RECT 441.530 498.400 441.670 499.160 ;
        RECT 441.530 498.200 441.990 498.400 ;
        RECT 441.670 498.140 441.990 498.200 ;
        RECT 441.670 472.840 441.990 472.900 ;
        RECT 441.300 472.700 441.990 472.840 ;
        RECT 441.300 471.820 441.440 472.700 ;
        RECT 441.670 472.640 441.990 472.700 ;
        RECT 442.590 471.820 442.910 471.880 ;
        RECT 441.300 471.680 442.910 471.820 ;
        RECT 442.590 471.620 442.910 471.680 ;
        RECT 442.590 16.900 442.910 16.960 ;
        RECT 463.290 16.900 463.610 16.960 ;
        RECT 442.590 16.760 463.610 16.900 ;
        RECT 442.590 16.700 442.910 16.760 ;
        RECT 463.290 16.700 463.610 16.760 ;
      LAYER via ;
        RECT 441.470 499.160 441.730 499.420 ;
        RECT 441.700 498.140 441.960 498.400 ;
        RECT 441.700 472.640 441.960 472.900 ;
        RECT 442.620 471.620 442.880 471.880 ;
        RECT 442.620 16.700 442.880 16.960 ;
        RECT 463.320 16.700 463.580 16.960 ;
      LAYER met2 ;
        RECT 441.490 500.000 441.770 504.000 ;
        RECT 441.530 499.450 441.670 500.000 ;
        RECT 441.470 499.130 441.730 499.450 ;
        RECT 441.700 498.110 441.960 498.430 ;
        RECT 441.760 472.930 441.900 498.110 ;
        RECT 441.700 472.610 441.960 472.930 ;
        RECT 442.620 471.590 442.880 471.910 ;
        RECT 442.680 16.990 442.820 471.590 ;
        RECT 442.620 16.670 442.880 16.990 ;
        RECT 463.320 16.670 463.580 16.990 ;
        RECT 463.380 2.400 463.520 16.670 ;
        RECT 463.170 -4.800 463.730 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.820 499.700 443.140 499.760 ;
        RECT 442.820 499.560 444.430 499.700 ;
        RECT 442.820 499.500 443.140 499.560 ;
        RECT 444.290 498.000 444.430 499.560 ;
        RECT 444.290 497.860 445.580 498.000 ;
        RECT 445.440 497.720 445.580 497.860 ;
        RECT 445.350 497.460 445.670 497.720 ;
        RECT 442.130 488.140 442.450 488.200 ;
        RECT 445.350 488.140 445.670 488.200 ;
        RECT 442.130 488.000 445.670 488.140 ;
        RECT 442.130 487.940 442.450 488.000 ;
        RECT 445.350 487.940 445.670 488.000 ;
        RECT 442.130 20.640 442.450 20.700 ;
        RECT 479.850 20.640 480.170 20.700 ;
        RECT 442.130 20.500 480.170 20.640 ;
        RECT 442.130 20.440 442.450 20.500 ;
        RECT 479.850 20.440 480.170 20.500 ;
      LAYER via ;
        RECT 442.850 499.500 443.110 499.760 ;
        RECT 445.380 497.460 445.640 497.720 ;
        RECT 442.160 487.940 442.420 488.200 ;
        RECT 445.380 487.940 445.640 488.200 ;
        RECT 442.160 20.440 442.420 20.700 ;
        RECT 479.880 20.440 480.140 20.700 ;
      LAYER met2 ;
        RECT 442.870 500.000 443.150 504.000 ;
        RECT 442.910 499.790 443.050 500.000 ;
        RECT 442.850 499.470 443.110 499.790 ;
        RECT 445.380 497.430 445.640 497.750 ;
        RECT 445.440 488.230 445.580 497.430 ;
        RECT 442.160 487.910 442.420 488.230 ;
        RECT 445.380 487.910 445.640 488.230 ;
        RECT 442.220 20.730 442.360 487.910 ;
        RECT 442.160 20.410 442.420 20.730 ;
        RECT 479.880 20.410 480.140 20.730 ;
        RECT 479.940 2.400 480.080 20.410 ;
        RECT 479.730 -4.800 480.290 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 416.600 499.360 416.920 499.420 ;
        RECT 416.600 499.220 417.750 499.360 ;
        RECT 416.600 499.160 416.920 499.220 ;
        RECT 417.610 498.400 417.750 499.220 ;
        RECT 417.610 498.200 418.070 498.400 ;
        RECT 417.750 498.140 418.070 498.200 ;
        RECT 417.750 472.160 418.070 472.220 ;
        RECT 418.670 472.160 418.990 472.220 ;
        RECT 417.750 472.020 418.990 472.160 ;
        RECT 417.750 471.960 418.070 472.020 ;
        RECT 418.670 471.960 418.990 472.020 ;
        RECT 378.650 20.640 378.970 20.700 ;
        RECT 418.670 20.640 418.990 20.700 ;
        RECT 378.650 20.500 418.990 20.640 ;
        RECT 378.650 20.440 378.970 20.500 ;
        RECT 418.670 20.440 418.990 20.500 ;
        RECT 165.210 17.920 165.530 17.980 ;
        RECT 378.650 17.920 378.970 17.980 ;
        RECT 165.210 17.780 378.970 17.920 ;
        RECT 165.210 17.720 165.530 17.780 ;
        RECT 378.650 17.720 378.970 17.780 ;
      LAYER via ;
        RECT 416.630 499.160 416.890 499.420 ;
        RECT 417.780 498.140 418.040 498.400 ;
        RECT 417.780 471.960 418.040 472.220 ;
        RECT 418.700 471.960 418.960 472.220 ;
        RECT 378.680 20.440 378.940 20.700 ;
        RECT 418.700 20.440 418.960 20.700 ;
        RECT 165.240 17.720 165.500 17.980 ;
        RECT 378.680 17.720 378.940 17.980 ;
      LAYER met2 ;
        RECT 416.650 500.000 416.930 504.000 ;
        RECT 416.690 499.450 416.830 500.000 ;
        RECT 416.630 499.130 416.890 499.450 ;
        RECT 417.780 498.110 418.040 498.430 ;
        RECT 417.840 472.250 417.980 498.110 ;
        RECT 417.780 471.930 418.040 472.250 ;
        RECT 418.700 471.930 418.960 472.250 ;
        RECT 418.760 20.730 418.900 471.930 ;
        RECT 378.680 20.410 378.940 20.730 ;
        RECT 418.700 20.410 418.960 20.730 ;
        RECT 378.740 18.010 378.880 20.410 ;
        RECT 165.240 17.690 165.500 18.010 ;
        RECT 378.680 17.690 378.940 18.010 ;
        RECT 165.300 2.400 165.440 17.690 ;
        RECT 165.090 -4.800 165.650 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.970 473.320 444.290 473.580 ;
        RECT 441.670 472.160 441.990 472.220 ;
        RECT 444.060 472.160 444.200 473.320 ;
        RECT 441.670 472.020 444.200 472.160 ;
        RECT 441.670 471.960 441.990 472.020 ;
        RECT 441.670 19.280 441.990 19.340 ;
        RECT 496.410 19.280 496.730 19.340 ;
        RECT 441.670 19.140 496.730 19.280 ;
        RECT 441.670 19.080 441.990 19.140 ;
        RECT 496.410 19.080 496.730 19.140 ;
      LAYER via ;
        RECT 444.000 473.320 444.260 473.580 ;
        RECT 441.700 471.960 441.960 472.220 ;
        RECT 441.700 19.080 441.960 19.340 ;
        RECT 496.440 19.080 496.700 19.340 ;
      LAYER met2 ;
        RECT 444.250 500.000 444.530 504.000 ;
        RECT 444.290 498.850 444.430 500.000 ;
        RECT 444.290 498.710 444.660 498.850 ;
        RECT 444.520 498.170 444.660 498.710 ;
        RECT 444.060 498.030 444.660 498.170 ;
        RECT 444.060 473.610 444.200 498.030 ;
        RECT 444.000 473.290 444.260 473.610 ;
        RECT 441.700 471.930 441.960 472.250 ;
        RECT 441.760 19.370 441.900 471.930 ;
        RECT 441.700 19.050 441.960 19.370 ;
        RECT 496.440 19.050 496.700 19.370 ;
        RECT 496.500 2.400 496.640 19.050 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 471.820 443.370 471.880 ;
        RECT 448.110 471.820 448.430 471.880 ;
        RECT 443.050 471.680 448.430 471.820 ;
        RECT 443.050 471.620 443.370 471.680 ;
        RECT 448.110 471.620 448.430 471.680 ;
        RECT 443.050 18.600 443.370 18.660 ;
        RECT 512.970 18.600 513.290 18.660 ;
        RECT 443.050 18.460 513.290 18.600 ;
        RECT 443.050 18.400 443.370 18.460 ;
        RECT 512.970 18.400 513.290 18.460 ;
      LAYER via ;
        RECT 443.080 471.620 443.340 471.880 ;
        RECT 448.140 471.620 448.400 471.880 ;
        RECT 443.080 18.400 443.340 18.660 ;
        RECT 513.000 18.400 513.260 18.660 ;
      LAYER met2 ;
        RECT 445.630 500.000 445.910 504.000 ;
        RECT 445.670 499.815 445.810 500.000 ;
        RECT 445.600 499.445 445.880 499.815 ;
        RECT 448.130 489.075 448.410 489.445 ;
        RECT 448.200 471.910 448.340 489.075 ;
        RECT 443.080 471.590 443.340 471.910 ;
        RECT 448.140 471.590 448.400 471.910 ;
        RECT 443.140 18.690 443.280 471.590 ;
        RECT 443.080 18.370 443.340 18.690 ;
        RECT 513.000 18.370 513.260 18.690 ;
        RECT 513.060 2.400 513.200 18.370 ;
        RECT 512.850 -4.800 513.410 2.400 ;
      LAYER via2 ;
        RECT 445.600 499.490 445.880 499.770 ;
        RECT 448.130 489.120 448.410 489.400 ;
      LAYER met3 ;
        RECT 445.575 499.620 445.905 499.795 ;
        RECT 445.550 499.610 445.930 499.620 ;
        RECT 445.550 499.310 446.190 499.610 ;
        RECT 445.550 499.300 445.930 499.310 ;
        RECT 445.550 489.410 445.930 489.420 ;
        RECT 448.105 489.410 448.435 489.425 ;
        RECT 445.550 489.110 448.435 489.410 ;
        RECT 445.550 489.100 445.930 489.110 ;
        RECT 448.105 489.095 448.435 489.110 ;
      LAYER via3 ;
        RECT 445.580 499.300 445.900 499.620 ;
        RECT 445.580 489.100 445.900 489.420 ;
      LAYER met4 ;
        RECT 445.575 499.295 445.905 499.625 ;
        RECT 445.590 489.425 445.890 499.295 ;
        RECT 445.575 489.095 445.905 489.425 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.010 500.000 447.290 504.000 ;
        RECT 447.050 499.020 447.190 500.000 ;
        RECT 446.820 498.880 447.190 499.020 ;
        RECT 446.820 498.285 446.960 498.880 ;
        RECT 446.750 497.915 447.030 498.285 ;
        RECT 529.550 17.155 529.830 17.525 ;
        RECT 529.620 2.400 529.760 17.155 ;
        RECT 529.410 -4.800 529.970 2.400 ;
      LAYER via2 ;
        RECT 446.750 497.960 447.030 498.240 ;
        RECT 529.550 17.200 529.830 17.480 ;
      LAYER met3 ;
        RECT 446.725 498.250 447.055 498.265 ;
        RECT 447.390 498.250 447.770 498.260 ;
        RECT 446.725 497.950 447.770 498.250 ;
        RECT 446.725 497.935 447.055 497.950 ;
        RECT 447.390 497.940 447.770 497.950 ;
        RECT 447.390 17.490 447.770 17.500 ;
        RECT 529.525 17.490 529.855 17.505 ;
        RECT 447.390 17.190 529.855 17.490 ;
        RECT 447.390 17.180 447.770 17.190 ;
        RECT 529.525 17.175 529.855 17.190 ;
      LAYER via3 ;
        RECT 447.420 497.940 447.740 498.260 ;
        RECT 447.420 17.180 447.740 17.500 ;
      LAYER met4 ;
        RECT 447.415 497.935 447.745 498.265 ;
        RECT 447.430 17.505 447.730 497.935 ;
        RECT 447.415 17.175 447.745 17.505 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 461.450 18.940 461.770 19.000 ;
        RECT 546.090 18.940 546.410 19.000 ;
        RECT 461.450 18.800 546.410 18.940 ;
        RECT 461.450 18.740 461.770 18.800 ;
        RECT 546.090 18.740 546.410 18.800 ;
      LAYER via ;
        RECT 461.480 18.740 461.740 19.000 ;
        RECT 546.120 18.740 546.380 19.000 ;
      LAYER met2 ;
        RECT 448.390 500.000 448.670 504.000 ;
        RECT 448.430 499.020 448.570 500.000 ;
        RECT 448.200 498.880 448.570 499.020 ;
        RECT 448.200 490.125 448.340 498.880 ;
        RECT 448.130 489.755 448.410 490.125 ;
        RECT 461.470 489.755 461.750 490.125 ;
        RECT 461.540 19.030 461.680 489.755 ;
        RECT 461.480 18.710 461.740 19.030 ;
        RECT 546.120 18.710 546.380 19.030 ;
        RECT 546.180 2.400 546.320 18.710 ;
        RECT 545.970 -4.800 546.530 2.400 ;
      LAYER via2 ;
        RECT 448.130 489.800 448.410 490.080 ;
        RECT 461.470 489.800 461.750 490.080 ;
      LAYER met3 ;
        RECT 448.105 490.090 448.435 490.105 ;
        RECT 461.445 490.090 461.775 490.105 ;
        RECT 448.105 489.790 461.775 490.090 ;
        RECT 448.105 489.775 448.435 489.790 ;
        RECT 461.445 489.775 461.775 489.790 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.950 488.480 450.270 488.540 ;
        RECT 455.470 488.480 455.790 488.540 ;
        RECT 449.950 488.340 455.790 488.480 ;
        RECT 449.950 488.280 450.270 488.340 ;
        RECT 455.470 488.280 455.790 488.340 ;
        RECT 455.470 472.160 455.790 472.220 ;
        RECT 459.610 472.160 459.930 472.220 ;
        RECT 455.470 472.020 459.930 472.160 ;
        RECT 455.470 471.960 455.790 472.020 ;
        RECT 459.610 471.960 459.930 472.020 ;
        RECT 459.610 17.920 459.930 17.980 ;
        RECT 562.650 17.920 562.970 17.980 ;
        RECT 459.610 17.780 562.970 17.920 ;
        RECT 459.610 17.720 459.930 17.780 ;
        RECT 562.650 17.720 562.970 17.780 ;
      LAYER via ;
        RECT 449.980 488.280 450.240 488.540 ;
        RECT 455.500 488.280 455.760 488.540 ;
        RECT 455.500 471.960 455.760 472.220 ;
        RECT 459.640 471.960 459.900 472.220 ;
        RECT 459.640 17.720 459.900 17.980 ;
        RECT 562.680 17.720 562.940 17.980 ;
      LAYER met2 ;
        RECT 449.770 500.000 450.050 504.000 ;
        RECT 449.810 498.340 449.950 500.000 ;
        RECT 449.810 498.200 450.180 498.340 ;
        RECT 450.040 488.570 450.180 498.200 ;
        RECT 449.980 488.250 450.240 488.570 ;
        RECT 455.500 488.250 455.760 488.570 ;
        RECT 455.560 472.250 455.700 488.250 ;
        RECT 455.500 471.930 455.760 472.250 ;
        RECT 459.640 471.930 459.900 472.250 ;
        RECT 459.700 18.010 459.840 471.930 ;
        RECT 459.640 17.690 459.900 18.010 ;
        RECT 562.680 17.690 562.940 18.010 ;
        RECT 562.740 2.400 562.880 17.690 ;
        RECT 562.530 -4.800 563.090 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.100 499.160 451.420 499.420 ;
        RECT 451.190 497.320 451.330 499.160 ;
        RECT 453.630 497.320 453.950 497.380 ;
        RECT 451.190 497.180 453.950 497.320 ;
        RECT 453.630 497.120 453.950 497.180 ;
        RECT 453.630 17.920 453.950 17.980 ;
        RECT 453.630 17.780 458.460 17.920 ;
        RECT 453.630 17.720 453.950 17.780 ;
        RECT 458.320 17.580 458.460 17.780 ;
        RECT 579.210 17.580 579.530 17.640 ;
        RECT 458.320 17.440 579.530 17.580 ;
        RECT 579.210 17.380 579.530 17.440 ;
      LAYER via ;
        RECT 451.130 499.160 451.390 499.420 ;
        RECT 453.660 497.120 453.920 497.380 ;
        RECT 453.660 17.720 453.920 17.980 ;
        RECT 579.240 17.380 579.500 17.640 ;
      LAYER met2 ;
        RECT 451.150 500.000 451.430 504.000 ;
        RECT 451.190 499.450 451.330 500.000 ;
        RECT 451.130 499.130 451.390 499.450 ;
        RECT 453.660 497.090 453.920 497.410 ;
        RECT 453.720 18.010 453.860 497.090 ;
        RECT 453.660 17.690 453.920 18.010 ;
        RECT 579.240 17.350 579.500 17.670 ;
        RECT 579.300 2.400 579.440 17.350 ;
        RECT 579.090 -4.800 579.650 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 452.480 500.380 452.800 500.440 ;
        RECT 450.730 500.240 452.800 500.380 ;
        RECT 450.730 496.980 450.870 500.240 ;
        RECT 452.480 500.180 452.800 500.240 ;
        RECT 454.090 496.980 454.410 497.040 ;
        RECT 450.730 496.840 454.410 496.980 ;
        RECT 454.090 496.780 454.410 496.840 ;
        RECT 454.090 487.120 454.410 487.180 ;
        RECT 460.070 487.120 460.390 487.180 ;
        RECT 454.090 486.980 460.390 487.120 ;
        RECT 454.090 486.920 454.410 486.980 ;
        RECT 460.070 486.920 460.390 486.980 ;
        RECT 460.070 24.380 460.390 24.440 ;
        RECT 595.770 24.380 596.090 24.440 ;
        RECT 460.070 24.240 596.090 24.380 ;
        RECT 460.070 24.180 460.390 24.240 ;
        RECT 595.770 24.180 596.090 24.240 ;
      LAYER via ;
        RECT 452.510 500.180 452.770 500.440 ;
        RECT 454.120 496.780 454.380 497.040 ;
        RECT 454.120 486.920 454.380 487.180 ;
        RECT 460.100 486.920 460.360 487.180 ;
        RECT 460.100 24.180 460.360 24.440 ;
        RECT 595.800 24.180 596.060 24.440 ;
      LAYER met2 ;
        RECT 452.530 500.470 452.810 504.000 ;
        RECT 452.510 500.150 452.810 500.470 ;
        RECT 452.530 500.000 452.810 500.150 ;
        RECT 454.120 496.750 454.380 497.070 ;
        RECT 454.180 487.210 454.320 496.750 ;
        RECT 454.120 486.890 454.380 487.210 ;
        RECT 460.100 486.890 460.360 487.210 ;
        RECT 460.160 24.470 460.300 486.890 ;
        RECT 460.100 24.150 460.360 24.470 ;
        RECT 595.800 24.150 596.060 24.470 ;
        RECT 595.860 2.400 596.000 24.150 ;
        RECT 595.650 -4.800 596.210 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.910 500.000 454.190 504.000 ;
        RECT 453.950 498.965 454.090 500.000 ;
        RECT 453.880 498.595 454.160 498.965 ;
        RECT 612.350 23.955 612.630 24.325 ;
        RECT 612.420 2.400 612.560 23.955 ;
        RECT 612.210 -4.800 612.770 2.400 ;
      LAYER via2 ;
        RECT 453.880 498.640 454.160 498.920 ;
        RECT 612.350 24.000 612.630 24.280 ;
      LAYER met3 ;
        RECT 453.855 498.940 454.185 498.945 ;
        RECT 453.830 498.930 454.210 498.940 ;
        RECT 453.400 498.630 454.210 498.930 ;
        RECT 453.830 498.620 454.210 498.630 ;
        RECT 453.855 498.615 454.185 498.620 ;
        RECT 453.830 24.290 454.210 24.300 ;
        RECT 612.325 24.290 612.655 24.305 ;
        RECT 453.830 23.990 612.655 24.290 ;
        RECT 453.830 23.980 454.210 23.990 ;
        RECT 612.325 23.975 612.655 23.990 ;
      LAYER via3 ;
        RECT 453.860 498.620 454.180 498.940 ;
        RECT 453.860 23.980 454.180 24.300 ;
      LAYER met4 ;
        RECT 453.855 498.615 454.185 498.945 ;
        RECT 453.870 24.305 454.170 498.615 ;
        RECT 453.855 23.975 454.185 24.305 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 489.500 455.790 489.560 ;
        RECT 460.530 489.500 460.850 489.560 ;
        RECT 455.470 489.360 460.850 489.500 ;
        RECT 455.470 489.300 455.790 489.360 ;
        RECT 460.530 489.300 460.850 489.360 ;
        RECT 460.530 18.260 460.850 18.320 ;
        RECT 628.890 18.260 629.210 18.320 ;
        RECT 460.530 18.120 629.210 18.260 ;
        RECT 460.530 18.060 460.850 18.120 ;
        RECT 628.890 18.060 629.210 18.120 ;
      LAYER via ;
        RECT 455.500 489.300 455.760 489.560 ;
        RECT 460.560 489.300 460.820 489.560 ;
        RECT 460.560 18.060 460.820 18.320 ;
        RECT 628.920 18.060 629.180 18.320 ;
      LAYER met2 ;
        RECT 455.290 500.000 455.570 504.000 ;
        RECT 455.330 498.680 455.470 500.000 ;
        RECT 455.330 498.540 455.700 498.680 ;
        RECT 455.560 489.590 455.700 498.540 ;
        RECT 455.500 489.270 455.760 489.590 ;
        RECT 460.560 489.270 460.820 489.590 ;
        RECT 460.620 18.350 460.760 489.270 ;
        RECT 460.560 18.030 460.820 18.350 ;
        RECT 628.920 18.030 629.180 18.350 ;
        RECT 628.980 2.400 629.120 18.030 ;
        RECT 628.770 -4.800 629.330 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.620 498.820 456.940 499.080 ;
        RECT 455.930 498.340 456.250 498.400 ;
        RECT 456.710 498.340 456.850 498.820 ;
        RECT 455.930 498.200 456.850 498.340 ;
        RECT 455.930 498.140 456.250 498.200 ;
        RECT 455.930 32.880 456.250 32.940 ;
        RECT 645.450 32.880 645.770 32.940 ;
        RECT 455.930 32.740 645.770 32.880 ;
        RECT 455.930 32.680 456.250 32.740 ;
        RECT 645.450 32.680 645.770 32.740 ;
      LAYER via ;
        RECT 456.650 498.820 456.910 499.080 ;
        RECT 455.960 498.140 456.220 498.400 ;
        RECT 455.960 32.680 456.220 32.940 ;
        RECT 645.480 32.680 645.740 32.940 ;
      LAYER met2 ;
        RECT 456.670 500.000 456.950 504.000 ;
        RECT 456.710 499.110 456.850 500.000 ;
        RECT 456.650 498.790 456.910 499.110 ;
        RECT 455.960 498.110 456.220 498.430 ;
        RECT 456.020 32.970 456.160 498.110 ;
        RECT 455.960 32.650 456.220 32.970 ;
        RECT 645.480 32.650 645.740 32.970 ;
        RECT 645.540 2.400 645.680 32.650 ;
        RECT 645.330 -4.800 645.890 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 415.450 472.840 415.770 472.900 ;
        RECT 417.290 472.840 417.610 472.900 ;
        RECT 415.450 472.700 417.610 472.840 ;
        RECT 415.450 472.640 415.770 472.700 ;
        RECT 417.290 472.640 417.610 472.700 ;
        RECT 187.290 18.260 187.610 18.320 ;
        RECT 415.450 18.260 415.770 18.320 ;
        RECT 187.290 18.120 415.770 18.260 ;
        RECT 187.290 18.060 187.610 18.120 ;
        RECT 415.450 18.060 415.770 18.120 ;
      LAYER via ;
        RECT 415.480 472.640 415.740 472.900 ;
        RECT 417.320 472.640 417.580 472.900 ;
        RECT 187.320 18.060 187.580 18.320 ;
        RECT 415.480 18.060 415.740 18.320 ;
      LAYER met2 ;
        RECT 418.490 500.000 418.770 504.000 ;
        RECT 418.530 499.645 418.670 500.000 ;
        RECT 418.460 499.275 418.740 499.645 ;
        RECT 417.310 496.615 417.590 496.985 ;
        RECT 417.380 472.930 417.520 496.615 ;
        RECT 415.480 472.610 415.740 472.930 ;
        RECT 417.320 472.610 417.580 472.930 ;
        RECT 415.540 18.350 415.680 472.610 ;
        RECT 187.320 18.030 187.580 18.350 ;
        RECT 415.480 18.030 415.740 18.350 ;
        RECT 187.380 2.400 187.520 18.030 ;
        RECT 187.170 -4.800 187.730 2.400 ;
      LAYER via2 ;
        RECT 418.460 499.320 418.740 499.600 ;
        RECT 417.310 496.660 417.590 496.940 ;
      LAYER met3 ;
        RECT 418.435 499.610 418.765 499.625 ;
        RECT 417.070 499.310 418.765 499.610 ;
        RECT 417.070 496.965 417.370 499.310 ;
        RECT 418.435 499.295 418.765 499.310 ;
        RECT 417.070 496.650 417.615 496.965 ;
        RECT 417.285 496.635 417.615 496.650 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.000 499.160 458.320 499.420 ;
        RECT 458.090 498.060 458.230 499.160 ;
        RECT 458.090 497.860 458.550 498.060 ;
        RECT 458.230 497.800 458.550 497.860 ;
        RECT 457.770 485.420 458.090 485.480 ;
        RECT 473.870 485.420 474.190 485.480 ;
        RECT 457.770 485.280 474.190 485.420 ;
        RECT 457.770 485.220 458.090 485.280 ;
        RECT 473.870 485.220 474.190 485.280 ;
        RECT 473.870 210.700 474.190 210.760 ;
        RECT 656.030 210.700 656.350 210.760 ;
        RECT 473.870 210.560 656.350 210.700 ;
        RECT 473.870 210.500 474.190 210.560 ;
        RECT 656.030 210.500 656.350 210.560 ;
        RECT 656.030 20.640 656.350 20.700 ;
        RECT 662.010 20.640 662.330 20.700 ;
        RECT 656.030 20.500 662.330 20.640 ;
        RECT 656.030 20.440 656.350 20.500 ;
        RECT 662.010 20.440 662.330 20.500 ;
      LAYER via ;
        RECT 458.030 499.160 458.290 499.420 ;
        RECT 458.260 497.800 458.520 498.060 ;
        RECT 457.800 485.220 458.060 485.480 ;
        RECT 473.900 485.220 474.160 485.480 ;
        RECT 473.900 210.500 474.160 210.760 ;
        RECT 656.060 210.500 656.320 210.760 ;
        RECT 656.060 20.440 656.320 20.700 ;
        RECT 662.040 20.440 662.300 20.700 ;
      LAYER met2 ;
        RECT 458.050 500.000 458.330 504.000 ;
        RECT 458.090 499.450 458.230 500.000 ;
        RECT 458.030 499.130 458.290 499.450 ;
        RECT 458.260 498.000 458.520 498.090 ;
        RECT 457.860 497.860 458.520 498.000 ;
        RECT 457.860 485.510 458.000 497.860 ;
        RECT 458.260 497.770 458.520 497.860 ;
        RECT 457.800 485.190 458.060 485.510 ;
        RECT 473.900 485.190 474.160 485.510 ;
        RECT 473.960 210.790 474.100 485.190 ;
        RECT 473.900 210.470 474.160 210.790 ;
        RECT 656.060 210.470 656.320 210.790 ;
        RECT 656.120 20.730 656.260 210.470 ;
        RECT 656.060 20.410 656.320 20.730 ;
        RECT 662.040 20.410 662.300 20.730 ;
        RECT 662.100 2.400 662.240 20.410 ;
        RECT 661.890 -4.800 662.450 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.850 473.180 457.170 473.240 ;
        RECT 459.150 473.180 459.470 473.240 ;
        RECT 456.850 473.040 459.470 473.180 ;
        RECT 456.850 472.980 457.170 473.040 ;
        RECT 459.150 472.980 459.470 473.040 ;
        RECT 456.850 438.160 457.170 438.220 ;
        RECT 576.910 438.160 577.230 438.220 ;
        RECT 456.850 438.020 577.230 438.160 ;
        RECT 456.850 437.960 457.170 438.020 ;
        RECT 576.910 437.960 577.230 438.020 ;
        RECT 576.910 19.620 577.230 19.680 ;
        RECT 678.570 19.620 678.890 19.680 ;
        RECT 576.910 19.480 678.890 19.620 ;
        RECT 576.910 19.420 577.230 19.480 ;
        RECT 678.570 19.420 678.890 19.480 ;
      LAYER via ;
        RECT 456.880 472.980 457.140 473.240 ;
        RECT 459.180 472.980 459.440 473.240 ;
        RECT 456.880 437.960 457.140 438.220 ;
        RECT 576.940 437.960 577.200 438.220 ;
        RECT 576.940 19.420 577.200 19.680 ;
        RECT 678.600 19.420 678.860 19.680 ;
      LAYER met2 ;
        RECT 459.430 500.000 459.710 504.000 ;
        RECT 459.470 499.815 459.610 500.000 ;
        RECT 459.400 499.445 459.680 499.815 ;
        RECT 459.170 498.595 459.450 498.965 ;
        RECT 459.240 473.270 459.380 498.595 ;
        RECT 456.880 472.950 457.140 473.270 ;
        RECT 459.180 472.950 459.440 473.270 ;
        RECT 456.940 438.250 457.080 472.950 ;
        RECT 456.880 437.930 457.140 438.250 ;
        RECT 576.940 437.930 577.200 438.250 ;
        RECT 577.000 19.710 577.140 437.930 ;
        RECT 576.940 19.390 577.200 19.710 ;
        RECT 678.600 19.390 678.860 19.710 ;
        RECT 678.660 2.400 678.800 19.390 ;
        RECT 678.450 -4.800 679.010 2.400 ;
      LAYER via2 ;
        RECT 459.400 499.490 459.680 499.770 ;
        RECT 459.170 498.640 459.450 498.920 ;
      LAYER met3 ;
        RECT 459.375 499.465 459.705 499.795 ;
        RECT 459.390 498.945 459.690 499.465 ;
        RECT 459.145 498.630 459.690 498.945 ;
        RECT 459.145 498.615 459.475 498.630 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.280 499.500 420.600 499.760 ;
        RECT 419.130 497.660 419.450 497.720 ;
        RECT 420.370 497.660 420.510 499.500 ;
        RECT 419.130 497.520 420.510 497.660 ;
        RECT 419.130 497.460 419.450 497.520 ;
        RECT 209.370 18.600 209.690 18.660 ;
        RECT 419.590 18.600 419.910 18.660 ;
        RECT 209.370 18.460 419.910 18.600 ;
        RECT 209.370 18.400 209.690 18.460 ;
        RECT 419.590 18.400 419.910 18.460 ;
      LAYER via ;
        RECT 420.310 499.500 420.570 499.760 ;
        RECT 419.160 497.460 419.420 497.720 ;
        RECT 209.400 18.400 209.660 18.660 ;
        RECT 419.620 18.400 419.880 18.660 ;
      LAYER met2 ;
        RECT 420.330 500.000 420.610 504.000 ;
        RECT 420.370 499.790 420.510 500.000 ;
        RECT 420.310 499.470 420.570 499.790 ;
        RECT 419.160 497.430 419.420 497.750 ;
        RECT 419.220 82.870 419.360 497.430 ;
        RECT 419.220 82.730 419.820 82.870 ;
        RECT 419.680 18.690 419.820 82.730 ;
        RECT 209.400 18.370 209.660 18.690 ;
        RECT 419.620 18.370 419.880 18.690 ;
        RECT 209.460 2.400 209.600 18.370 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.170 500.000 422.450 504.000 ;
        RECT 422.210 499.645 422.350 500.000 ;
        RECT 422.140 499.275 422.420 499.645 ;
        RECT 231.470 23.955 231.750 24.325 ;
        RECT 231.540 2.400 231.680 23.955 ;
        RECT 231.330 -4.800 231.890 2.400 ;
      LAYER via2 ;
        RECT 422.140 499.320 422.420 499.600 ;
        RECT 231.470 24.000 231.750 24.280 ;
      LAYER met3 ;
        RECT 420.710 499.610 421.090 499.620 ;
        RECT 422.115 499.610 422.445 499.625 ;
        RECT 420.710 499.310 422.445 499.610 ;
        RECT 420.710 499.300 421.090 499.310 ;
        RECT 422.115 499.295 422.445 499.310 ;
        RECT 231.445 24.290 231.775 24.305 ;
        RECT 419.790 24.290 420.170 24.300 ;
        RECT 231.445 23.990 420.170 24.290 ;
        RECT 231.445 23.975 231.775 23.990 ;
        RECT 419.790 23.980 420.170 23.990 ;
      LAYER via3 ;
        RECT 420.740 499.300 421.060 499.620 ;
        RECT 419.820 23.980 420.140 24.300 ;
      LAYER met4 ;
        RECT 420.735 499.295 421.065 499.625 ;
        RECT 420.750 448.650 421.050 499.295 ;
        RECT 419.830 448.350 421.050 448.650 ;
        RECT 419.830 24.305 420.130 448.350 ;
        RECT 419.815 23.975 420.145 24.305 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.500 499.160 423.820 499.420 ;
        RECT 422.350 497.660 422.670 497.720 ;
        RECT 423.590 497.660 423.730 499.160 ;
        RECT 422.350 497.520 423.730 497.660 ;
        RECT 422.350 497.460 422.670 497.520 ;
        RECT 248.010 25.060 248.330 25.120 ;
        RECT 422.350 25.060 422.670 25.120 ;
        RECT 248.010 24.920 422.670 25.060 ;
        RECT 248.010 24.860 248.330 24.920 ;
        RECT 422.350 24.860 422.670 24.920 ;
      LAYER via ;
        RECT 423.530 499.160 423.790 499.420 ;
        RECT 422.380 497.460 422.640 497.720 ;
        RECT 248.040 24.860 248.300 25.120 ;
        RECT 422.380 24.860 422.640 25.120 ;
      LAYER met2 ;
        RECT 423.550 500.000 423.830 504.000 ;
        RECT 423.590 499.450 423.730 500.000 ;
        RECT 423.530 499.130 423.790 499.450 ;
        RECT 422.380 497.430 422.640 497.750 ;
        RECT 422.440 25.150 422.580 497.430 ;
        RECT 248.040 24.830 248.300 25.150 ;
        RECT 422.380 24.830 422.640 25.150 ;
        RECT 248.100 2.400 248.240 24.830 ;
        RECT 247.890 -4.800 248.450 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 425.110 473.520 425.430 473.580 ;
        RECT 426.950 473.520 427.270 473.580 ;
        RECT 425.110 473.380 427.270 473.520 ;
        RECT 425.110 473.320 425.430 473.380 ;
        RECT 426.950 473.320 427.270 473.380 ;
        RECT 264.570 25.740 264.890 25.800 ;
        RECT 426.950 25.740 427.270 25.800 ;
        RECT 264.570 25.600 427.270 25.740 ;
        RECT 264.570 25.540 264.890 25.600 ;
        RECT 426.950 25.540 427.270 25.600 ;
      LAYER via ;
        RECT 425.140 473.320 425.400 473.580 ;
        RECT 426.980 473.320 427.240 473.580 ;
        RECT 264.600 25.540 264.860 25.800 ;
        RECT 426.980 25.540 427.240 25.800 ;
      LAYER met2 ;
        RECT 424.930 500.000 425.210 504.000 ;
        RECT 424.970 498.340 425.110 500.000 ;
        RECT 424.970 498.200 425.340 498.340 ;
        RECT 425.200 473.610 425.340 498.200 ;
        RECT 425.140 473.290 425.400 473.610 ;
        RECT 426.980 473.290 427.240 473.610 ;
        RECT 427.040 25.830 427.180 473.290 ;
        RECT 264.600 25.510 264.860 25.830 ;
        RECT 426.980 25.510 427.240 25.830 ;
        RECT 264.660 2.400 264.800 25.510 ;
        RECT 264.450 -4.800 265.010 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.650 497.320 424.970 497.380 ;
        RECT 426.030 497.320 426.350 497.380 ;
        RECT 424.650 497.180 426.350 497.320 ;
        RECT 424.650 497.120 424.970 497.180 ;
        RECT 426.030 497.120 426.350 497.180 ;
        RECT 281.130 26.080 281.450 26.140 ;
        RECT 425.110 26.080 425.430 26.140 ;
        RECT 281.130 25.940 425.430 26.080 ;
        RECT 281.130 25.880 281.450 25.940 ;
        RECT 425.110 25.880 425.430 25.940 ;
      LAYER via ;
        RECT 424.680 497.120 424.940 497.380 ;
        RECT 426.060 497.120 426.320 497.380 ;
        RECT 281.160 25.880 281.420 26.140 ;
        RECT 425.140 25.880 425.400 26.140 ;
      LAYER met2 ;
        RECT 426.310 500.000 426.590 504.000 ;
        RECT 426.350 498.850 426.490 500.000 ;
        RECT 426.120 498.710 426.490 498.850 ;
        RECT 426.120 497.410 426.260 498.710 ;
        RECT 424.680 497.090 424.940 497.410 ;
        RECT 426.060 497.090 426.320 497.410 ;
        RECT 424.740 472.840 424.880 497.090 ;
        RECT 424.740 472.700 425.340 472.840 ;
        RECT 425.200 26.170 425.340 472.700 ;
        RECT 281.160 25.850 281.420 26.170 ;
        RECT 425.140 25.850 425.400 26.170 ;
        RECT 281.220 2.400 281.360 25.850 ;
        RECT 281.010 -4.800 281.570 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.690 500.000 427.970 504.000 ;
        RECT 427.730 499.645 427.870 500.000 ;
        RECT 427.660 499.275 427.940 499.645 ;
        RECT 297.710 24.635 297.990 25.005 ;
        RECT 297.780 2.400 297.920 24.635 ;
        RECT 297.570 -4.800 298.130 2.400 ;
      LAYER via2 ;
        RECT 427.660 499.320 427.940 499.600 ;
        RECT 297.710 24.680 297.990 24.960 ;
      LAYER met3 ;
        RECT 427.635 499.610 427.965 499.625 ;
        RECT 427.635 499.295 428.180 499.610 ;
        RECT 427.880 498.940 428.180 499.295 ;
        RECT 427.880 498.630 428.450 498.940 ;
        RECT 428.070 498.620 428.450 498.630 ;
        RECT 297.685 24.970 298.015 24.985 ;
        RECT 428.070 24.970 428.450 24.980 ;
        RECT 297.685 24.670 428.450 24.970 ;
        RECT 297.685 24.655 298.015 24.670 ;
        RECT 428.070 24.660 428.450 24.670 ;
      LAYER via3 ;
        RECT 428.100 498.620 428.420 498.940 ;
        RECT 428.100 24.660 428.420 24.980 ;
      LAYER met4 ;
        RECT 428.095 498.615 428.425 498.945 ;
        RECT 428.110 24.985 428.410 498.615 ;
        RECT 428.095 24.655 428.425 24.985 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.020 499.160 429.340 499.420 ;
        RECT 426.490 498.000 426.810 498.060 ;
        RECT 429.110 498.000 429.250 499.160 ;
        RECT 426.490 497.860 429.250 498.000 ;
        RECT 426.490 497.800 426.810 497.860 ;
        RECT 424.190 472.160 424.510 472.220 ;
        RECT 426.490 472.160 426.810 472.220 ;
        RECT 424.190 472.020 426.810 472.160 ;
        RECT 424.190 471.960 424.510 472.020 ;
        RECT 426.490 471.960 426.810 472.020 ;
        RECT 314.250 32.200 314.570 32.260 ;
        RECT 424.190 32.200 424.510 32.260 ;
        RECT 314.250 32.060 424.510 32.200 ;
        RECT 314.250 32.000 314.570 32.060 ;
        RECT 424.190 32.000 424.510 32.060 ;
      LAYER via ;
        RECT 429.050 499.160 429.310 499.420 ;
        RECT 426.520 497.800 426.780 498.060 ;
        RECT 424.220 471.960 424.480 472.220 ;
        RECT 426.520 471.960 426.780 472.220 ;
        RECT 314.280 32.000 314.540 32.260 ;
        RECT 424.220 32.000 424.480 32.260 ;
      LAYER met2 ;
        RECT 429.070 500.000 429.350 504.000 ;
        RECT 429.110 499.450 429.250 500.000 ;
        RECT 429.050 499.130 429.310 499.450 ;
        RECT 426.520 497.770 426.780 498.090 ;
        RECT 426.580 472.250 426.720 497.770 ;
        RECT 424.220 471.930 424.480 472.250 ;
        RECT 426.520 471.930 426.780 472.250 ;
        RECT 424.280 32.290 424.420 471.930 ;
        RECT 314.280 31.970 314.540 32.290 ;
        RECT 424.220 31.970 424.480 32.290 ;
        RECT 314.340 2.400 314.480 31.970 ;
        RECT 314.130 -4.800 314.690 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 126.570 24.720 126.890 24.780 ;
        RECT 412.230 24.720 412.550 24.780 ;
        RECT 126.570 24.580 412.550 24.720 ;
        RECT 126.570 24.520 126.890 24.580 ;
        RECT 412.230 24.520 412.550 24.580 ;
      LAYER via ;
        RECT 126.600 24.520 126.860 24.780 ;
        RECT 412.260 24.520 412.520 24.780 ;
      LAYER met2 ;
        RECT 413.430 500.000 413.710 504.000 ;
        RECT 413.470 498.850 413.610 500.000 ;
        RECT 413.240 498.710 413.610 498.850 ;
        RECT 413.240 496.870 413.380 498.710 ;
        RECT 412.780 496.730 413.380 496.870 ;
        RECT 412.780 472.840 412.920 496.730 ;
        RECT 412.320 472.700 412.920 472.840 ;
        RECT 412.320 24.810 412.460 472.700 ;
        RECT 126.600 24.490 126.860 24.810 ;
        RECT 412.260 24.490 412.520 24.810 ;
        RECT 126.660 2.400 126.800 24.490 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 415.220 499.160 415.540 499.420 ;
        RECT 415.310 498.340 415.450 499.160 ;
        RECT 415.910 498.340 416.230 498.400 ;
        RECT 415.310 498.200 416.230 498.340 ;
        RECT 415.910 498.140 416.230 498.200 ;
        RECT 400.270 26.420 400.590 26.480 ;
        RECT 415.910 26.420 416.230 26.480 ;
        RECT 400.270 26.280 416.230 26.420 ;
        RECT 400.270 26.220 400.590 26.280 ;
        RECT 415.910 26.220 416.230 26.280 ;
        RECT 400.270 17.920 400.590 17.980 ;
        RECT 379.200 17.780 400.590 17.920 ;
        RECT 379.200 17.580 379.340 17.780 ;
        RECT 400.270 17.720 400.590 17.780 ;
        RECT 161.620 17.440 379.340 17.580 ;
        RECT 148.650 17.240 148.970 17.300 ;
        RECT 161.620 17.240 161.760 17.440 ;
        RECT 148.650 17.100 161.760 17.240 ;
        RECT 148.650 17.040 148.970 17.100 ;
      LAYER via ;
        RECT 415.250 499.160 415.510 499.420 ;
        RECT 415.940 498.140 416.200 498.400 ;
        RECT 400.300 26.220 400.560 26.480 ;
        RECT 415.940 26.220 416.200 26.480 ;
        RECT 400.300 17.720 400.560 17.980 ;
        RECT 148.680 17.040 148.940 17.300 ;
      LAYER met2 ;
        RECT 415.270 500.000 415.550 504.000 ;
        RECT 415.310 499.450 415.450 500.000 ;
        RECT 415.250 499.130 415.510 499.450 ;
        RECT 415.940 498.110 416.200 498.430 ;
        RECT 416.000 26.510 416.140 498.110 ;
        RECT 400.300 26.190 400.560 26.510 ;
        RECT 415.940 26.190 416.200 26.510 ;
        RECT 400.360 18.010 400.500 26.190 ;
        RECT 400.300 17.690 400.560 18.010 ;
        RECT 148.680 17.010 148.940 17.330 ;
        RECT 148.740 2.400 148.880 17.010 ;
        RECT 148.530 -4.800 149.090 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.860 499.500 431.180 499.760 ;
        RECT 430.950 497.040 431.090 499.500 ;
        RECT 430.950 496.840 431.410 497.040 ;
        RECT 431.090 496.780 431.410 496.840 ;
        RECT 336.330 32.880 336.650 32.940 ;
        RECT 431.090 32.880 431.410 32.940 ;
        RECT 336.330 32.740 431.410 32.880 ;
        RECT 336.330 32.680 336.650 32.740 ;
        RECT 431.090 32.680 431.410 32.740 ;
      LAYER via ;
        RECT 430.890 499.500 431.150 499.760 ;
        RECT 431.120 496.780 431.380 497.040 ;
        RECT 336.360 32.680 336.620 32.940 ;
        RECT 431.120 32.680 431.380 32.940 ;
      LAYER met2 ;
        RECT 430.910 500.000 431.190 504.000 ;
        RECT 430.950 499.790 431.090 500.000 ;
        RECT 430.890 499.470 431.150 499.790 ;
        RECT 431.120 496.750 431.380 497.070 ;
        RECT 431.180 32.970 431.320 496.750 ;
        RECT 336.360 32.650 336.620 32.970 ;
        RECT 431.120 32.650 431.380 32.970 ;
        RECT 336.420 2.400 336.560 32.650 ;
        RECT 336.210 -4.800 336.770 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.240 498.820 432.560 499.080 ;
        RECT 432.330 498.060 432.470 498.820 ;
        RECT 432.010 497.860 432.470 498.060 ;
        RECT 432.010 497.800 432.330 497.860 ;
        RECT 421.890 487.120 422.210 487.180 ;
        RECT 432.010 487.120 432.330 487.180 ;
        RECT 421.890 486.980 432.330 487.120 ;
        RECT 421.890 486.920 422.210 486.980 ;
        RECT 432.010 486.920 432.330 486.980 ;
        RECT 421.890 471.820 422.210 471.880 ;
        RECT 424.650 471.820 424.970 471.880 ;
        RECT 421.890 471.680 424.970 471.820 ;
        RECT 421.890 471.620 422.210 471.680 ;
        RECT 424.650 471.620 424.970 471.680 ;
        RECT 352.890 33.560 353.210 33.620 ;
        RECT 424.650 33.560 424.970 33.620 ;
        RECT 352.890 33.420 424.970 33.560 ;
        RECT 352.890 33.360 353.210 33.420 ;
        RECT 424.650 33.360 424.970 33.420 ;
      LAYER via ;
        RECT 432.270 498.820 432.530 499.080 ;
        RECT 432.040 497.800 432.300 498.060 ;
        RECT 421.920 486.920 422.180 487.180 ;
        RECT 432.040 486.920 432.300 487.180 ;
        RECT 421.920 471.620 422.180 471.880 ;
        RECT 424.680 471.620 424.940 471.880 ;
        RECT 352.920 33.360 353.180 33.620 ;
        RECT 424.680 33.360 424.940 33.620 ;
      LAYER met2 ;
        RECT 432.290 500.000 432.570 504.000 ;
        RECT 432.330 499.110 432.470 500.000 ;
        RECT 432.270 498.790 432.530 499.110 ;
        RECT 432.040 497.770 432.300 498.090 ;
        RECT 432.100 487.210 432.240 497.770 ;
        RECT 421.920 486.890 422.180 487.210 ;
        RECT 432.040 486.890 432.300 487.210 ;
        RECT 421.980 471.910 422.120 486.890 ;
        RECT 421.920 471.590 422.180 471.910 ;
        RECT 424.680 471.590 424.940 471.910 ;
        RECT 424.740 33.650 424.880 471.590 ;
        RECT 352.920 33.330 353.180 33.650 ;
        RECT 424.680 33.330 424.940 33.650 ;
        RECT 352.980 2.400 353.120 33.330 ;
        RECT 352.770 -4.800 353.330 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 433.620 499.020 433.940 499.080 ;
        RECT 433.620 498.820 434.080 499.020 ;
        RECT 433.940 498.400 434.080 498.820 ;
        RECT 433.850 498.140 434.170 498.400 ;
        RECT 429.710 471.820 430.030 471.880 ;
        RECT 433.850 471.820 434.170 471.880 ;
        RECT 429.710 471.680 434.170 471.820 ;
        RECT 429.710 471.620 430.030 471.680 ;
        RECT 433.850 471.620 434.170 471.680 ;
        RECT 369.450 33.900 369.770 33.960 ;
        RECT 429.710 33.900 430.030 33.960 ;
        RECT 369.450 33.760 430.030 33.900 ;
        RECT 369.450 33.700 369.770 33.760 ;
        RECT 429.710 33.700 430.030 33.760 ;
      LAYER via ;
        RECT 433.650 498.820 433.910 499.080 ;
        RECT 433.880 498.140 434.140 498.400 ;
        RECT 429.740 471.620 430.000 471.880 ;
        RECT 433.880 471.620 434.140 471.880 ;
        RECT 369.480 33.700 369.740 33.960 ;
        RECT 429.740 33.700 430.000 33.960 ;
      LAYER met2 ;
        RECT 433.670 500.000 433.950 504.000 ;
        RECT 433.710 499.110 433.850 500.000 ;
        RECT 433.650 498.790 433.910 499.110 ;
        RECT 433.880 498.110 434.140 498.430 ;
        RECT 433.940 471.910 434.080 498.110 ;
        RECT 429.740 471.590 430.000 471.910 ;
        RECT 433.880 471.590 434.140 471.910 ;
        RECT 429.800 33.990 429.940 471.590 ;
        RECT 369.480 33.670 369.740 33.990 ;
        RECT 429.740 33.670 430.000 33.990 ;
        RECT 369.540 2.400 369.680 33.670 ;
        RECT 369.330 -4.800 369.890 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.000 499.500 435.320 499.760 ;
        RECT 435.090 497.660 435.230 499.500 ;
        RECT 437.070 497.660 437.390 497.720 ;
        RECT 435.090 497.520 437.390 497.660 ;
        RECT 437.070 497.460 437.390 497.520 ;
        RECT 437.070 483.720 437.390 483.780 ;
        RECT 431.180 483.580 437.390 483.720 ;
        RECT 428.330 483.040 428.650 483.100 ;
        RECT 431.180 483.040 431.320 483.580 ;
        RECT 437.070 483.520 437.390 483.580 ;
        RECT 428.330 482.900 431.320 483.040 ;
        RECT 428.330 482.840 428.650 482.900 ;
        RECT 379.570 417.420 379.890 417.480 ;
        RECT 427.870 417.420 428.190 417.480 ;
        RECT 379.570 417.280 428.190 417.420 ;
        RECT 379.570 417.220 379.890 417.280 ;
        RECT 427.870 417.220 428.190 417.280 ;
        RECT 379.570 17.580 379.890 17.640 ;
        RECT 386.010 17.580 386.330 17.640 ;
        RECT 379.570 17.440 386.330 17.580 ;
        RECT 379.570 17.380 379.890 17.440 ;
        RECT 386.010 17.380 386.330 17.440 ;
      LAYER via ;
        RECT 435.030 499.500 435.290 499.760 ;
        RECT 437.100 497.460 437.360 497.720 ;
        RECT 428.360 482.840 428.620 483.100 ;
        RECT 437.100 483.520 437.360 483.780 ;
        RECT 379.600 417.220 379.860 417.480 ;
        RECT 427.900 417.220 428.160 417.480 ;
        RECT 379.600 17.380 379.860 17.640 ;
        RECT 386.040 17.380 386.300 17.640 ;
      LAYER met2 ;
        RECT 435.050 500.000 435.330 504.000 ;
        RECT 435.090 499.790 435.230 500.000 ;
        RECT 435.030 499.470 435.290 499.790 ;
        RECT 437.100 497.430 437.360 497.750 ;
        RECT 437.160 483.810 437.300 497.430 ;
        RECT 437.100 483.490 437.360 483.810 ;
        RECT 428.360 482.810 428.620 483.130 ;
        RECT 428.420 420.970 428.560 482.810 ;
        RECT 427.960 420.830 428.560 420.970 ;
        RECT 427.960 417.510 428.100 420.830 ;
        RECT 379.600 417.190 379.860 417.510 ;
        RECT 427.900 417.190 428.160 417.510 ;
        RECT 379.660 17.670 379.800 417.190 ;
        RECT 379.600 17.350 379.860 17.670 ;
        RECT 386.040 17.350 386.300 17.670 ;
        RECT 386.100 2.400 386.240 17.350 ;
        RECT 385.890 -4.800 386.450 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.380 498.820 436.700 499.080 ;
        RECT 436.470 498.000 436.610 498.820 ;
        RECT 436.470 497.860 438.220 498.000 ;
        RECT 438.080 497.720 438.220 497.860 ;
        RECT 437.990 497.460 438.310 497.720 ;
        RECT 411.770 24.040 412.090 24.100 ;
        RECT 438.450 24.040 438.770 24.100 ;
        RECT 411.770 23.900 438.770 24.040 ;
        RECT 411.770 23.840 412.090 23.900 ;
        RECT 438.450 23.840 438.770 23.900 ;
        RECT 402.570 14.180 402.890 14.240 ;
        RECT 411.770 14.180 412.090 14.240 ;
        RECT 402.570 14.040 412.090 14.180 ;
        RECT 402.570 13.980 402.890 14.040 ;
        RECT 411.770 13.980 412.090 14.040 ;
      LAYER via ;
        RECT 436.410 498.820 436.670 499.080 ;
        RECT 438.020 497.460 438.280 497.720 ;
        RECT 411.800 23.840 412.060 24.100 ;
        RECT 438.480 23.840 438.740 24.100 ;
        RECT 402.600 13.980 402.860 14.240 ;
        RECT 411.800 13.980 412.060 14.240 ;
      LAYER met2 ;
        RECT 436.430 500.000 436.710 504.000 ;
        RECT 436.470 499.110 436.610 500.000 ;
        RECT 436.410 498.790 436.670 499.110 ;
        RECT 438.020 497.430 438.280 497.750 ;
        RECT 438.080 473.690 438.220 497.430 ;
        RECT 438.080 473.550 438.680 473.690 ;
        RECT 438.540 24.130 438.680 473.550 ;
        RECT 411.800 23.810 412.060 24.130 ;
        RECT 438.480 23.810 438.740 24.130 ;
        RECT 411.860 14.270 412.000 23.810 ;
        RECT 402.600 13.950 402.860 14.270 ;
        RECT 411.800 13.950 412.060 14.270 ;
        RECT 402.660 2.400 402.800 13.950 ;
        RECT 402.450 -4.800 403.010 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 437.760 499.160 438.080 499.420 ;
        RECT 437.850 499.020 437.990 499.160 ;
        RECT 437.620 498.880 437.990 499.020 ;
        RECT 437.620 498.740 437.760 498.880 ;
        RECT 437.530 498.480 437.850 498.740 ;
        RECT 432.010 483.380 432.330 483.440 ;
        RECT 437.530 483.380 437.850 483.440 ;
        RECT 432.010 483.240 437.850 483.380 ;
        RECT 432.010 483.180 432.330 483.240 ;
        RECT 437.530 483.180 437.850 483.240 ;
        RECT 417.750 421.160 418.070 421.220 ;
        RECT 432.010 421.160 432.330 421.220 ;
        RECT 417.750 421.020 432.330 421.160 ;
        RECT 417.750 420.960 418.070 421.020 ;
        RECT 432.010 420.960 432.330 421.020 ;
      LAYER via ;
        RECT 437.790 499.160 438.050 499.420 ;
        RECT 437.560 498.480 437.820 498.740 ;
        RECT 432.040 483.180 432.300 483.440 ;
        RECT 437.560 483.180 437.820 483.440 ;
        RECT 417.780 420.960 418.040 421.220 ;
        RECT 432.040 420.960 432.300 421.220 ;
      LAYER met2 ;
        RECT 437.810 500.000 438.090 504.000 ;
        RECT 437.850 499.450 437.990 500.000 ;
        RECT 437.790 499.130 438.050 499.450 ;
        RECT 437.560 498.450 437.820 498.770 ;
        RECT 437.620 483.470 437.760 498.450 ;
        RECT 432.040 483.150 432.300 483.470 ;
        RECT 437.560 483.150 437.820 483.470 ;
        RECT 432.100 421.250 432.240 483.150 ;
        RECT 417.780 420.930 418.040 421.250 ;
        RECT 432.040 420.930 432.300 421.250 ;
        RECT 417.840 82.870 417.980 420.930 ;
        RECT 417.840 82.730 418.440 82.870 ;
        RECT 418.300 17.410 418.440 82.730 ;
        RECT 418.300 17.270 419.360 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 439.140 499.500 439.460 499.760 ;
        RECT 439.230 498.400 439.370 499.500 ;
        RECT 439.230 498.200 439.690 498.400 ;
        RECT 439.370 498.140 439.690 498.200 ;
      LAYER via ;
        RECT 439.170 499.500 439.430 499.760 ;
        RECT 439.400 498.140 439.660 498.400 ;
      LAYER met2 ;
        RECT 439.190 500.000 439.470 504.000 ;
        RECT 439.230 499.790 439.370 500.000 ;
        RECT 439.170 499.470 439.430 499.790 ;
        RECT 439.400 498.340 439.660 498.430 ;
        RECT 439.400 498.200 440.060 498.340 ;
        RECT 439.400 498.110 439.660 498.200 ;
        RECT 439.920 34.570 440.060 498.200 ;
        RECT 439.000 34.430 440.060 34.570 ;
        RECT 439.000 2.450 439.140 34.430 ;
        RECT 435.570 1.770 436.130 2.400 ;
        RECT 438.080 2.310 439.140 2.450 ;
        RECT 438.080 1.770 438.220 2.310 ;
        RECT 435.570 1.630 438.220 1.770 ;
        RECT 435.570 -4.800 436.130 1.630 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 437.070 472.500 437.390 472.560 ;
        RECT 440.290 472.500 440.610 472.560 ;
        RECT 437.070 472.360 440.610 472.500 ;
        RECT 437.070 472.300 437.390 472.360 ;
        RECT 440.290 472.300 440.610 472.360 ;
        RECT 437.070 17.240 437.390 17.300 ;
        RECT 452.250 17.240 452.570 17.300 ;
        RECT 437.070 17.100 452.570 17.240 ;
        RECT 437.070 17.040 437.390 17.100 ;
        RECT 452.250 17.040 452.570 17.100 ;
      LAYER via ;
        RECT 437.100 472.300 437.360 472.560 ;
        RECT 440.320 472.300 440.580 472.560 ;
        RECT 437.100 17.040 437.360 17.300 ;
        RECT 452.280 17.040 452.540 17.300 ;
      LAYER met2 ;
        RECT 440.570 500.000 440.850 504.000 ;
        RECT 440.610 499.645 440.750 500.000 ;
        RECT 440.540 499.275 440.820 499.645 ;
        RECT 440.310 497.915 440.590 498.285 ;
        RECT 440.380 472.590 440.520 497.915 ;
        RECT 437.100 472.270 437.360 472.590 ;
        RECT 440.320 472.270 440.580 472.590 ;
        RECT 437.160 17.330 437.300 472.270 ;
        RECT 437.100 17.010 437.360 17.330 ;
        RECT 452.280 17.010 452.540 17.330 ;
        RECT 452.340 2.400 452.480 17.010 ;
        RECT 452.130 -4.800 452.690 2.400 ;
      LAYER via2 ;
        RECT 440.540 499.320 440.820 499.600 ;
        RECT 440.310 497.960 440.590 498.240 ;
      LAYER met3 ;
        RECT 440.515 499.610 440.845 499.625 ;
        RECT 439.610 499.310 440.845 499.610 ;
        RECT 439.610 498.250 439.910 499.310 ;
        RECT 440.515 499.295 440.845 499.310 ;
        RECT 440.285 498.250 440.615 498.265 ;
        RECT 439.610 497.950 440.615 498.250 ;
        RECT 440.285 497.935 440.615 497.950 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.970 20.980 444.290 21.040 ;
        RECT 468.810 20.980 469.130 21.040 ;
        RECT 443.970 20.840 469.130 20.980 ;
        RECT 443.970 20.780 444.290 20.840 ;
        RECT 468.810 20.780 469.130 20.840 ;
      LAYER via ;
        RECT 444.000 20.780 444.260 21.040 ;
        RECT 468.840 20.780 469.100 21.040 ;
      LAYER met2 ;
        RECT 441.950 500.000 442.230 504.000 ;
        RECT 441.990 499.135 442.130 500.000 ;
        RECT 441.920 498.765 442.200 499.135 ;
        RECT 442.610 497.235 442.890 497.605 ;
        RECT 442.680 491.880 442.820 497.235 ;
        RECT 442.680 491.740 443.280 491.880 ;
        RECT 443.140 473.010 443.280 491.740 ;
        RECT 443.140 472.870 444.200 473.010 ;
        RECT 444.060 21.070 444.200 472.870 ;
        RECT 444.000 20.750 444.260 21.070 ;
        RECT 468.840 20.750 469.100 21.070 ;
        RECT 468.900 2.400 469.040 20.750 ;
        RECT 468.690 -4.800 469.250 2.400 ;
      LAYER via2 ;
        RECT 441.920 498.810 442.200 499.090 ;
        RECT 442.610 497.280 442.890 497.560 ;
      LAYER met3 ;
        RECT 441.895 498.785 442.225 499.115 ;
        RECT 441.910 497.570 442.210 498.785 ;
        RECT 442.585 497.570 442.915 497.585 ;
        RECT 441.910 497.270 442.915 497.570 ;
        RECT 442.585 497.255 442.915 497.270 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 492.560 443.370 492.620 ;
        RECT 444.430 492.560 444.750 492.620 ;
        RECT 443.050 492.420 444.750 492.560 ;
        RECT 443.050 492.360 443.370 492.420 ;
        RECT 444.430 492.360 444.750 492.420 ;
        RECT 444.430 26.420 444.750 26.480 ;
        RECT 485.370 26.420 485.690 26.480 ;
        RECT 444.430 26.280 485.690 26.420 ;
        RECT 444.430 26.220 444.750 26.280 ;
        RECT 485.370 26.220 485.690 26.280 ;
      LAYER via ;
        RECT 443.080 492.360 443.340 492.620 ;
        RECT 444.460 492.360 444.720 492.620 ;
        RECT 444.460 26.220 444.720 26.480 ;
        RECT 485.400 26.220 485.660 26.480 ;
      LAYER met2 ;
        RECT 443.330 500.000 443.610 504.000 ;
        RECT 443.370 498.680 443.510 500.000 ;
        RECT 443.140 498.540 443.510 498.680 ;
        RECT 443.140 492.650 443.280 498.540 ;
        RECT 443.080 492.330 443.340 492.650 ;
        RECT 444.460 492.330 444.720 492.650 ;
        RECT 444.520 26.510 444.660 492.330 ;
        RECT 444.460 26.190 444.720 26.510 ;
        RECT 485.400 26.190 485.660 26.510 ;
        RECT 485.460 2.400 485.600 26.190 ;
        RECT 485.250 -4.800 485.810 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 170.730 30.840 171.050 30.900 ;
        RECT 416.370 30.840 416.690 30.900 ;
        RECT 170.730 30.700 416.690 30.840 ;
        RECT 170.730 30.640 171.050 30.700 ;
        RECT 416.370 30.640 416.690 30.700 ;
      LAYER via ;
        RECT 170.760 30.640 171.020 30.900 ;
        RECT 416.400 30.640 416.660 30.900 ;
      LAYER met2 ;
        RECT 417.110 500.000 417.390 504.000 ;
        RECT 417.150 498.850 417.290 500.000 ;
        RECT 416.920 498.710 417.290 498.850 ;
        RECT 416.920 498.170 417.060 498.710 ;
        RECT 416.460 498.030 417.060 498.170 ;
        RECT 416.460 30.930 416.600 498.030 ;
        RECT 170.760 30.610 171.020 30.930 ;
        RECT 416.400 30.610 416.660 30.930 ;
        RECT 170.820 2.400 170.960 30.610 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.660 499.700 444.980 499.760 ;
        RECT 444.660 499.500 445.120 499.700 ;
        RECT 444.980 498.400 445.120 499.500 ;
        RECT 444.890 498.140 445.210 498.400 ;
        RECT 444.890 27.440 445.210 27.500 ;
        RECT 501.930 27.440 502.250 27.500 ;
        RECT 444.890 27.300 502.250 27.440 ;
        RECT 444.890 27.240 445.210 27.300 ;
        RECT 501.930 27.240 502.250 27.300 ;
      LAYER via ;
        RECT 444.690 499.500 444.950 499.760 ;
        RECT 444.920 498.140 445.180 498.400 ;
        RECT 444.920 27.240 445.180 27.500 ;
        RECT 501.960 27.240 502.220 27.500 ;
      LAYER met2 ;
        RECT 444.710 500.000 444.990 504.000 ;
        RECT 444.750 499.790 444.890 500.000 ;
        RECT 444.690 499.470 444.950 499.790 ;
        RECT 444.920 498.110 445.180 498.430 ;
        RECT 444.980 27.530 445.120 498.110 ;
        RECT 444.920 27.210 445.180 27.530 ;
        RECT 501.960 27.210 502.220 27.530 ;
        RECT 502.020 2.400 502.160 27.210 ;
        RECT 501.810 -4.800 502.370 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.040 499.500 446.360 499.760 ;
        RECT 446.130 498.740 446.270 499.500 ;
        RECT 445.810 498.540 446.270 498.740 ;
        RECT 445.810 498.480 446.130 498.540 ;
        RECT 446.270 491.880 446.590 491.940 ;
        RECT 454.550 491.880 454.870 491.940 ;
        RECT 446.270 491.740 454.870 491.880 ;
        RECT 446.270 491.680 446.590 491.740 ;
        RECT 454.550 491.680 454.870 491.740 ;
        RECT 454.090 26.760 454.410 26.820 ;
        RECT 454.090 26.620 494.340 26.760 ;
        RECT 454.090 26.560 454.410 26.620 ;
        RECT 494.200 26.080 494.340 26.620 ;
        RECT 518.490 26.080 518.810 26.140 ;
        RECT 494.200 25.940 518.810 26.080 ;
        RECT 518.490 25.880 518.810 25.940 ;
      LAYER via ;
        RECT 446.070 499.500 446.330 499.760 ;
        RECT 445.840 498.480 446.100 498.740 ;
        RECT 446.300 491.680 446.560 491.940 ;
        RECT 454.580 491.680 454.840 491.940 ;
        RECT 454.120 26.560 454.380 26.820 ;
        RECT 518.520 25.880 518.780 26.140 ;
      LAYER met2 ;
        RECT 446.090 500.000 446.370 504.000 ;
        RECT 446.130 499.790 446.270 500.000 ;
        RECT 446.070 499.470 446.330 499.790 ;
        RECT 445.840 498.680 446.100 498.770 ;
        RECT 445.840 498.540 446.500 498.680 ;
        RECT 445.840 498.450 446.100 498.540 ;
        RECT 446.360 491.970 446.500 498.540 ;
        RECT 446.300 491.650 446.560 491.970 ;
        RECT 454.580 491.650 454.840 491.970 ;
        RECT 454.640 420.970 454.780 491.650 ;
        RECT 454.180 420.830 454.780 420.970 ;
        RECT 454.180 26.850 454.320 420.830 ;
        RECT 454.120 26.530 454.380 26.850 ;
        RECT 518.520 25.850 518.780 26.170 ;
        RECT 518.580 2.400 518.720 25.850 ;
        RECT 518.370 -4.800 518.930 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 447.420 498.820 447.740 499.080 ;
        RECT 447.510 498.680 447.650 498.820 ;
        RECT 447.280 498.540 447.650 498.680 ;
        RECT 447.280 498.400 447.420 498.540 ;
        RECT 447.190 498.140 447.510 498.400 ;
        RECT 447.190 490.860 447.510 490.920 ;
        RECT 448.570 490.860 448.890 490.920 ;
        RECT 447.190 490.720 448.890 490.860 ;
        RECT 447.190 490.660 447.510 490.720 ;
        RECT 448.570 490.660 448.890 490.720 ;
        RECT 448.570 26.080 448.890 26.140 ;
        RECT 448.570 25.940 493.420 26.080 ;
        RECT 448.570 25.880 448.890 25.940 ;
        RECT 493.280 25.740 493.420 25.940 ;
        RECT 493.280 25.600 493.880 25.740 ;
        RECT 493.740 25.400 493.880 25.600 ;
        RECT 535.050 25.400 535.370 25.460 ;
        RECT 493.740 25.260 535.370 25.400 ;
        RECT 535.050 25.200 535.370 25.260 ;
      LAYER via ;
        RECT 447.450 498.820 447.710 499.080 ;
        RECT 447.220 498.140 447.480 498.400 ;
        RECT 447.220 490.660 447.480 490.920 ;
        RECT 448.600 490.660 448.860 490.920 ;
        RECT 448.600 25.880 448.860 26.140 ;
        RECT 535.080 25.200 535.340 25.460 ;
      LAYER met2 ;
        RECT 447.470 500.000 447.750 504.000 ;
        RECT 447.510 499.110 447.650 500.000 ;
        RECT 447.450 498.790 447.710 499.110 ;
        RECT 447.220 498.110 447.480 498.430 ;
        RECT 447.280 490.950 447.420 498.110 ;
        RECT 447.220 490.630 447.480 490.950 ;
        RECT 448.600 490.630 448.860 490.950 ;
        RECT 448.660 26.170 448.800 490.630 ;
        RECT 448.600 25.850 448.860 26.170 ;
        RECT 535.080 25.170 535.340 25.490 ;
        RECT 535.140 2.400 535.280 25.170 ;
        RECT 534.930 -4.800 535.490 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 491.540 448.890 491.600 ;
        RECT 449.490 491.540 449.810 491.600 ;
        RECT 448.570 491.400 449.810 491.540 ;
        RECT 448.570 491.340 448.890 491.400 ;
        RECT 449.490 491.340 449.810 491.400 ;
        RECT 449.950 25.400 450.270 25.460 ;
        RECT 449.950 25.260 478.240 25.400 ;
        RECT 449.950 25.200 450.270 25.260 ;
        RECT 478.100 24.720 478.240 25.260 ;
        RECT 551.610 24.720 551.930 24.780 ;
        RECT 478.100 24.580 551.930 24.720 ;
        RECT 551.610 24.520 551.930 24.580 ;
      LAYER via ;
        RECT 448.600 491.340 448.860 491.600 ;
        RECT 449.520 491.340 449.780 491.600 ;
        RECT 449.980 25.200 450.240 25.460 ;
        RECT 551.640 24.520 551.900 24.780 ;
      LAYER met2 ;
        RECT 448.850 500.000 449.130 504.000 ;
        RECT 448.890 498.680 449.030 500.000 ;
        RECT 448.660 498.540 449.030 498.680 ;
        RECT 448.660 491.630 448.800 498.540 ;
        RECT 448.600 491.310 448.860 491.630 ;
        RECT 449.520 491.310 449.780 491.630 ;
        RECT 449.580 473.010 449.720 491.310 ;
        RECT 449.580 472.870 450.180 473.010 ;
        RECT 450.040 25.490 450.180 472.870 ;
        RECT 449.980 25.170 450.240 25.490 ;
        RECT 551.640 24.490 551.900 24.810 ;
        RECT 551.700 2.400 551.840 24.490 ;
        RECT 551.490 -4.800 552.050 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.870 31.180 451.190 31.240 ;
        RECT 568.170 31.180 568.490 31.240 ;
        RECT 450.870 31.040 568.490 31.180 ;
        RECT 450.870 30.980 451.190 31.040 ;
        RECT 568.170 30.980 568.490 31.040 ;
      LAYER via ;
        RECT 450.900 30.980 451.160 31.240 ;
        RECT 568.200 30.980 568.460 31.240 ;
      LAYER met2 ;
        RECT 450.230 500.000 450.510 504.000 ;
        RECT 450.270 499.645 450.410 500.000 ;
        RECT 450.200 499.275 450.480 499.645 ;
        RECT 450.890 491.115 451.170 491.485 ;
        RECT 450.960 31.270 451.100 491.115 ;
        RECT 450.900 30.950 451.160 31.270 ;
        RECT 568.200 30.950 568.460 31.270 ;
        RECT 568.260 2.400 568.400 30.950 ;
        RECT 568.050 -4.800 568.610 2.400 ;
      LAYER via2 ;
        RECT 450.200 499.320 450.480 499.600 ;
        RECT 450.890 491.160 451.170 491.440 ;
      LAYER met3 ;
        RECT 450.175 499.620 450.505 499.625 ;
        RECT 450.150 499.610 450.530 499.620 ;
        RECT 450.150 499.310 450.960 499.610 ;
        RECT 450.150 499.300 450.530 499.310 ;
        RECT 450.175 499.295 450.505 499.300 ;
        RECT 450.150 491.450 450.530 491.460 ;
        RECT 450.865 491.450 451.195 491.465 ;
        RECT 450.150 491.150 451.195 491.450 ;
        RECT 450.150 491.140 450.530 491.150 ;
        RECT 450.865 491.135 451.195 491.150 ;
      LAYER via3 ;
        RECT 450.180 499.300 450.500 499.620 ;
        RECT 450.180 491.140 450.500 491.460 ;
      LAYER met4 ;
        RECT 450.175 499.295 450.505 499.625 ;
        RECT 450.190 491.465 450.490 499.295 ;
        RECT 450.175 491.135 450.505 491.465 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.560 499.500 451.880 499.760 ;
        RECT 451.650 498.740 451.790 499.500 ;
        RECT 451.650 498.540 452.110 498.740 ;
        RECT 451.790 498.480 452.110 498.540 ;
        RECT 450.410 472.840 450.730 472.900 ;
        RECT 451.330 472.840 451.650 472.900 ;
        RECT 450.410 472.700 451.650 472.840 ;
        RECT 450.410 472.640 450.730 472.700 ;
        RECT 451.330 472.640 451.650 472.700 ;
        RECT 450.410 30.840 450.730 30.900 ;
        RECT 584.730 30.840 585.050 30.900 ;
        RECT 450.410 30.700 585.050 30.840 ;
        RECT 450.410 30.640 450.730 30.700 ;
        RECT 584.730 30.640 585.050 30.700 ;
      LAYER via ;
        RECT 451.590 499.500 451.850 499.760 ;
        RECT 451.820 498.480 452.080 498.740 ;
        RECT 450.440 472.640 450.700 472.900 ;
        RECT 451.360 472.640 451.620 472.900 ;
        RECT 450.440 30.640 450.700 30.900 ;
        RECT 584.760 30.640 585.020 30.900 ;
      LAYER met2 ;
        RECT 451.610 500.000 451.890 504.000 ;
        RECT 451.650 499.790 451.790 500.000 ;
        RECT 451.590 499.470 451.850 499.790 ;
        RECT 451.820 498.680 452.080 498.770 ;
        RECT 451.420 498.540 452.080 498.680 ;
        RECT 451.420 472.930 451.560 498.540 ;
        RECT 451.820 498.450 452.080 498.540 ;
        RECT 450.440 472.610 450.700 472.930 ;
        RECT 451.360 472.610 451.620 472.930 ;
        RECT 450.500 30.930 450.640 472.610 ;
        RECT 450.440 30.610 450.700 30.930 ;
        RECT 584.760 30.610 585.020 30.930 ;
        RECT 584.820 2.400 584.960 30.610 ;
        RECT 584.610 -4.800 585.170 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 452.940 499.700 453.260 499.760 ;
        RECT 452.940 499.500 453.400 499.700 ;
        RECT 453.260 499.080 453.400 499.500 ;
        RECT 453.170 498.820 453.490 499.080 ;
        RECT 449.490 472.500 449.810 472.560 ;
        RECT 453.170 472.500 453.490 472.560 ;
        RECT 449.490 472.360 453.490 472.500 ;
        RECT 449.490 472.300 449.810 472.360 ;
        RECT 453.170 472.300 453.490 472.360 ;
        RECT 449.490 24.040 449.810 24.100 ;
        RECT 601.290 24.040 601.610 24.100 ;
        RECT 449.490 23.900 601.610 24.040 ;
        RECT 449.490 23.840 449.810 23.900 ;
        RECT 601.290 23.840 601.610 23.900 ;
      LAYER via ;
        RECT 452.970 499.500 453.230 499.760 ;
        RECT 453.200 498.820 453.460 499.080 ;
        RECT 449.520 472.300 449.780 472.560 ;
        RECT 453.200 472.300 453.460 472.560 ;
        RECT 449.520 23.840 449.780 24.100 ;
        RECT 601.320 23.840 601.580 24.100 ;
      LAYER met2 ;
        RECT 452.990 500.000 453.270 504.000 ;
        RECT 453.030 499.790 453.170 500.000 ;
        RECT 452.970 499.470 453.230 499.790 ;
        RECT 453.200 498.790 453.460 499.110 ;
        RECT 453.260 472.590 453.400 498.790 ;
        RECT 449.520 472.270 449.780 472.590 ;
        RECT 453.200 472.270 453.460 472.590 ;
        RECT 449.580 24.130 449.720 472.270 ;
        RECT 449.520 23.810 449.780 24.130 ;
        RECT 601.320 23.810 601.580 24.130 ;
        RECT 601.380 2.400 601.520 23.810 ;
        RECT 601.170 -4.800 601.730 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.170 18.600 522.490 18.660 ;
        RECT 617.850 18.600 618.170 18.660 ;
        RECT 522.170 18.460 618.170 18.600 ;
        RECT 522.170 18.400 522.490 18.460 ;
        RECT 617.850 18.400 618.170 18.460 ;
      LAYER via ;
        RECT 522.200 18.400 522.460 18.660 ;
        RECT 617.880 18.400 618.140 18.660 ;
      LAYER met2 ;
        RECT 454.370 500.000 454.650 504.000 ;
        RECT 453.650 498.170 453.930 498.285 ;
        RECT 454.410 498.170 454.550 500.000 ;
        RECT 453.650 498.030 454.550 498.170 ;
        RECT 453.650 497.915 453.930 498.030 ;
        RECT 522.190 437.395 522.470 437.765 ;
        RECT 522.260 18.690 522.400 437.395 ;
        RECT 522.200 18.370 522.460 18.690 ;
        RECT 617.880 18.370 618.140 18.690 ;
        RECT 617.940 2.400 618.080 18.370 ;
        RECT 617.730 -4.800 618.290 2.400 ;
      LAYER via2 ;
        RECT 453.650 497.960 453.930 498.240 ;
        RECT 522.190 437.440 522.470 437.720 ;
      LAYER met3 ;
        RECT 452.910 498.250 453.290 498.260 ;
        RECT 453.625 498.250 453.955 498.265 ;
        RECT 452.910 497.950 453.955 498.250 ;
        RECT 452.910 497.940 453.290 497.950 ;
        RECT 453.625 497.935 453.955 497.950 ;
        RECT 452.910 437.730 453.290 437.740 ;
        RECT 522.165 437.730 522.495 437.745 ;
        RECT 452.910 437.430 522.495 437.730 ;
        RECT 452.910 437.420 453.290 437.430 ;
        RECT 522.165 437.415 522.495 437.430 ;
      LAYER via3 ;
        RECT 452.940 497.940 453.260 498.260 ;
        RECT 452.940 437.420 453.260 437.740 ;
      LAYER met4 ;
        RECT 452.935 497.935 453.265 498.265 ;
        RECT 452.950 437.745 453.250 497.935 ;
        RECT 452.935 437.415 453.265 437.745 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.310 451.760 457.630 451.820 ;
        RECT 596.690 451.760 597.010 451.820 ;
        RECT 457.310 451.620 597.010 451.760 ;
        RECT 457.310 451.560 457.630 451.620 ;
        RECT 596.690 451.560 597.010 451.620 ;
        RECT 596.690 18.940 597.010 19.000 ;
        RECT 634.410 18.940 634.730 19.000 ;
        RECT 596.690 18.800 634.730 18.940 ;
        RECT 596.690 18.740 597.010 18.800 ;
        RECT 634.410 18.740 634.730 18.800 ;
      LAYER via ;
        RECT 457.340 451.560 457.600 451.820 ;
        RECT 596.720 451.560 596.980 451.820 ;
        RECT 596.720 18.740 596.980 19.000 ;
        RECT 634.440 18.740 634.700 19.000 ;
      LAYER met2 ;
        RECT 455.750 500.000 456.030 504.000 ;
        RECT 455.790 499.020 455.930 500.000 ;
        RECT 455.790 498.965 456.160 499.020 ;
        RECT 455.790 498.880 456.230 498.965 ;
        RECT 455.950 498.595 456.230 498.880 ;
        RECT 456.870 497.915 457.150 498.285 ;
        RECT 456.940 476.170 457.080 497.915 ;
        RECT 456.940 476.030 457.540 476.170 ;
        RECT 457.400 451.850 457.540 476.030 ;
        RECT 457.340 451.530 457.600 451.850 ;
        RECT 596.720 451.530 596.980 451.850 ;
        RECT 596.780 19.030 596.920 451.530 ;
        RECT 596.720 18.710 596.980 19.030 ;
        RECT 634.440 18.710 634.700 19.030 ;
        RECT 634.500 2.400 634.640 18.710 ;
        RECT 634.290 -4.800 634.850 2.400 ;
      LAYER via2 ;
        RECT 455.950 498.640 456.230 498.920 ;
        RECT 456.870 497.960 457.150 498.240 ;
      LAYER met3 ;
        RECT 455.925 498.930 456.255 498.945 ;
        RECT 455.710 498.615 456.255 498.930 ;
        RECT 455.710 498.250 456.010 498.615 ;
        RECT 456.845 498.250 457.175 498.265 ;
        RECT 455.710 497.950 457.175 498.250 ;
        RECT 456.845 497.935 457.175 497.950 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.310 490.860 457.630 490.920 ;
        RECT 457.310 490.720 463.980 490.860 ;
        RECT 457.310 490.660 457.630 490.720 ;
        RECT 463.840 489.840 463.980 490.720 ;
        RECT 463.840 489.700 545.170 489.840 ;
        RECT 545.030 489.500 545.170 489.700 ;
        RECT 648.670 489.500 648.990 489.560 ;
        RECT 545.030 489.360 648.990 489.500 ;
        RECT 648.670 489.300 648.990 489.360 ;
      LAYER via ;
        RECT 457.340 490.660 457.600 490.920 ;
        RECT 648.700 489.300 648.960 489.560 ;
      LAYER met2 ;
        RECT 457.130 500.000 457.410 504.000 ;
        RECT 457.170 498.680 457.310 500.000 ;
        RECT 457.170 498.540 457.540 498.680 ;
        RECT 457.400 490.950 457.540 498.540 ;
        RECT 457.340 490.630 457.600 490.950 ;
        RECT 648.700 489.270 648.960 489.590 ;
        RECT 648.760 82.870 648.900 489.270 ;
        RECT 648.760 82.730 651.200 82.870 ;
        RECT 651.060 2.400 651.200 82.730 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 418.900 498.820 419.220 499.080 ;
        RECT 418.210 498.340 418.530 498.400 ;
        RECT 418.990 498.340 419.130 498.820 ;
        RECT 418.210 498.200 419.130 498.340 ;
        RECT 418.210 498.140 418.530 498.200 ;
        RECT 416.830 473.520 417.150 473.580 ;
        RECT 418.210 473.520 418.530 473.580 ;
        RECT 416.830 473.380 418.530 473.520 ;
        RECT 416.830 473.320 417.150 473.380 ;
        RECT 418.210 473.320 418.530 473.380 ;
        RECT 192.810 31.180 193.130 31.240 ;
        RECT 416.830 31.180 417.150 31.240 ;
        RECT 192.810 31.040 417.150 31.180 ;
        RECT 192.810 30.980 193.130 31.040 ;
        RECT 416.830 30.980 417.150 31.040 ;
      LAYER via ;
        RECT 418.930 498.820 419.190 499.080 ;
        RECT 418.240 498.140 418.500 498.400 ;
        RECT 416.860 473.320 417.120 473.580 ;
        RECT 418.240 473.320 418.500 473.580 ;
        RECT 192.840 30.980 193.100 31.240 ;
        RECT 416.860 30.980 417.120 31.240 ;
      LAYER met2 ;
        RECT 418.950 500.000 419.230 504.000 ;
        RECT 418.990 499.110 419.130 500.000 ;
        RECT 418.930 498.790 419.190 499.110 ;
        RECT 418.240 498.110 418.500 498.430 ;
        RECT 418.300 473.610 418.440 498.110 ;
        RECT 416.860 473.290 417.120 473.610 ;
        RECT 418.240 473.290 418.500 473.610 ;
        RECT 416.920 31.270 417.060 473.290 ;
        RECT 192.840 30.950 193.100 31.270 ;
        RECT 416.860 30.950 417.120 31.270 ;
        RECT 192.900 2.400 193.040 30.950 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.790 488.820 659.110 488.880 ;
        RECT 467.290 488.680 659.110 488.820 ;
        RECT 458.230 488.480 458.550 488.540 ;
        RECT 467.290 488.480 467.430 488.680 ;
        RECT 658.790 488.620 659.110 488.680 ;
        RECT 458.230 488.340 467.430 488.480 ;
        RECT 458.230 488.280 458.550 488.340 ;
        RECT 658.790 16.220 659.110 16.280 ;
        RECT 667.530 16.220 667.850 16.280 ;
        RECT 658.790 16.080 667.850 16.220 ;
        RECT 658.790 16.020 659.110 16.080 ;
        RECT 667.530 16.020 667.850 16.080 ;
      LAYER via ;
        RECT 458.260 488.280 458.520 488.540 ;
        RECT 658.820 488.620 659.080 488.880 ;
        RECT 658.820 16.020 659.080 16.280 ;
        RECT 667.560 16.020 667.820 16.280 ;
      LAYER met2 ;
        RECT 458.510 500.000 458.790 504.000 ;
        RECT 458.550 498.680 458.690 500.000 ;
        RECT 458.550 498.540 458.920 498.680 ;
        RECT 458.780 491.200 458.920 498.540 ;
        RECT 458.320 491.060 458.920 491.200 ;
        RECT 458.320 488.570 458.460 491.060 ;
        RECT 658.820 488.590 659.080 488.910 ;
        RECT 458.260 488.250 458.520 488.570 ;
        RECT 658.880 16.310 659.020 488.590 ;
        RECT 658.820 15.990 659.080 16.310 ;
        RECT 667.560 15.990 667.820 16.310 ;
        RECT 667.620 2.400 667.760 15.990 ;
        RECT 667.410 -4.800 667.970 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 472.840 456.710 472.900 ;
        RECT 459.610 472.840 459.930 472.900 ;
        RECT 456.390 472.700 459.930 472.840 ;
        RECT 456.390 472.640 456.710 472.700 ;
        RECT 459.610 472.640 459.930 472.700 ;
        RECT 456.390 210.360 456.710 210.420 ;
        RECT 683.630 210.360 683.950 210.420 ;
        RECT 456.390 210.220 683.950 210.360 ;
        RECT 456.390 210.160 456.710 210.220 ;
        RECT 683.630 210.160 683.950 210.220 ;
      LAYER via ;
        RECT 456.420 472.640 456.680 472.900 ;
        RECT 459.640 472.640 459.900 472.900 ;
        RECT 456.420 210.160 456.680 210.420 ;
        RECT 683.660 210.160 683.920 210.420 ;
      LAYER met2 ;
        RECT 459.890 500.000 460.170 504.000 ;
        RECT 459.930 498.680 460.070 500.000 ;
        RECT 459.700 498.540 460.070 498.680 ;
        RECT 459.700 472.930 459.840 498.540 ;
        RECT 456.420 472.610 456.680 472.930 ;
        RECT 459.640 472.610 459.900 472.930 ;
        RECT 456.480 210.450 456.620 472.610 ;
        RECT 456.420 210.130 456.680 210.450 ;
        RECT 683.660 210.130 683.920 210.450 ;
        RECT 683.720 82.870 683.860 210.130 ;
        RECT 683.720 82.730 684.320 82.870 ;
        RECT 684.180 2.400 684.320 82.730 ;
        RECT 683.970 -4.800 684.530 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.740 499.500 421.060 499.760 ;
        RECT 420.830 498.740 420.970 499.500 ;
        RECT 420.830 498.540 421.290 498.740 ;
        RECT 420.970 498.480 421.290 498.540 ;
      LAYER via ;
        RECT 420.770 499.500 421.030 499.760 ;
        RECT 421.000 498.480 421.260 498.740 ;
      LAYER met2 ;
        RECT 420.790 500.000 421.070 504.000 ;
        RECT 420.830 499.790 420.970 500.000 ;
        RECT 420.770 499.470 421.030 499.790 ;
        RECT 421.000 498.450 421.260 498.770 ;
        RECT 421.060 491.485 421.200 498.450 ;
        RECT 420.990 491.115 421.270 491.485 ;
        RECT 214.910 37.555 215.190 37.925 ;
        RECT 214.980 2.400 215.120 37.555 ;
        RECT 214.770 -4.800 215.330 2.400 ;
      LAYER via2 ;
        RECT 420.990 491.160 421.270 491.440 ;
        RECT 214.910 37.600 215.190 37.880 ;
      LAYER met3 ;
        RECT 420.965 491.450 421.295 491.465 ;
        RECT 421.630 491.450 422.010 491.460 ;
        RECT 420.965 491.150 422.010 491.450 ;
        RECT 420.965 491.135 421.295 491.150 ;
        RECT 421.630 491.140 422.010 491.150 ;
        RECT 214.885 37.890 215.215 37.905 ;
        RECT 421.630 37.890 422.010 37.900 ;
        RECT 214.885 37.590 422.010 37.890 ;
        RECT 214.885 37.575 215.215 37.590 ;
        RECT 421.630 37.580 422.010 37.590 ;
      LAYER via3 ;
        RECT 421.660 491.140 421.980 491.460 ;
        RECT 421.660 37.580 421.980 37.900 ;
      LAYER met4 ;
        RECT 421.655 491.135 421.985 491.465 ;
        RECT 421.670 37.905 421.970 491.135 ;
        RECT 421.655 37.575 421.985 37.905 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 422.350 498.340 422.670 498.400 ;
        RECT 421.520 498.200 422.670 498.340 ;
        RECT 421.520 496.980 421.660 498.200 ;
        RECT 422.350 498.140 422.670 498.200 ;
        RECT 424.190 496.980 424.510 497.040 ;
        RECT 421.520 496.840 424.510 496.980 ;
        RECT 424.190 496.780 424.510 496.840 ;
        RECT 234.670 224.640 234.990 224.700 ;
        RECT 423.730 224.640 424.050 224.700 ;
        RECT 234.670 224.500 424.050 224.640 ;
        RECT 234.670 224.440 234.990 224.500 ;
        RECT 423.730 224.440 424.050 224.500 ;
      LAYER via ;
        RECT 422.380 498.140 422.640 498.400 ;
        RECT 424.220 496.780 424.480 497.040 ;
        RECT 234.700 224.440 234.960 224.700 ;
        RECT 423.760 224.440 424.020 224.700 ;
      LAYER met2 ;
        RECT 422.630 500.000 422.910 504.000 ;
        RECT 422.670 498.850 422.810 500.000 ;
        RECT 422.440 498.710 422.810 498.850 ;
        RECT 422.440 498.430 422.580 498.710 ;
        RECT 422.380 498.110 422.640 498.430 ;
        RECT 424.220 496.750 424.480 497.070 ;
        RECT 424.280 472.840 424.420 496.750 ;
        RECT 423.820 472.700 424.420 472.840 ;
        RECT 423.820 224.730 423.960 472.700 ;
        RECT 234.700 224.410 234.960 224.730 ;
        RECT 423.760 224.410 424.020 224.730 ;
        RECT 234.760 82.870 234.900 224.410 ;
        RECT 234.760 82.730 237.200 82.870 ;
        RECT 237.060 2.400 237.200 82.730 ;
        RECT 236.850 -4.800 237.410 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.730 473.860 424.050 473.920 ;
        RECT 425.570 473.860 425.890 473.920 ;
        RECT 423.730 473.720 425.890 473.860 ;
        RECT 423.730 473.660 424.050 473.720 ;
        RECT 425.570 473.660 425.890 473.720 ;
        RECT 253.530 25.400 253.850 25.460 ;
        RECT 425.570 25.400 425.890 25.460 ;
        RECT 253.530 25.260 425.890 25.400 ;
        RECT 253.530 25.200 253.850 25.260 ;
        RECT 425.570 25.200 425.890 25.260 ;
      LAYER via ;
        RECT 423.760 473.660 424.020 473.920 ;
        RECT 425.600 473.660 425.860 473.920 ;
        RECT 253.560 25.200 253.820 25.460 ;
        RECT 425.600 25.200 425.860 25.460 ;
      LAYER met2 ;
        RECT 424.010 500.000 424.290 504.000 ;
        RECT 424.050 498.850 424.190 500.000 ;
        RECT 423.820 498.710 424.190 498.850 ;
        RECT 423.820 473.950 423.960 498.710 ;
        RECT 423.760 473.630 424.020 473.950 ;
        RECT 425.600 473.630 425.860 473.950 ;
        RECT 425.660 25.490 425.800 473.630 ;
        RECT 253.560 25.170 253.820 25.490 ;
        RECT 425.600 25.170 425.860 25.490 ;
        RECT 253.620 2.400 253.760 25.170 ;
        RECT 253.410 -4.800 253.970 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.170 431.360 269.490 431.420 ;
        RECT 426.030 431.360 426.350 431.420 ;
        RECT 269.170 431.220 426.350 431.360 ;
        RECT 269.170 431.160 269.490 431.220 ;
        RECT 426.030 431.160 426.350 431.220 ;
      LAYER via ;
        RECT 269.200 431.160 269.460 431.420 ;
        RECT 426.060 431.160 426.320 431.420 ;
      LAYER met2 ;
        RECT 425.390 500.000 425.670 504.000 ;
        RECT 425.430 499.645 425.570 500.000 ;
        RECT 425.360 499.275 425.640 499.645 ;
        RECT 426.050 496.555 426.330 496.925 ;
        RECT 426.120 431.450 426.260 496.555 ;
        RECT 269.200 431.130 269.460 431.450 ;
        RECT 426.060 431.130 426.320 431.450 ;
        RECT 269.260 82.870 269.400 431.130 ;
        RECT 269.260 82.730 270.320 82.870 ;
        RECT 270.180 2.400 270.320 82.730 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 425.360 499.320 425.640 499.600 ;
        RECT 426.050 496.600 426.330 496.880 ;
      LAYER met3 ;
        RECT 425.335 499.620 425.665 499.625 ;
        RECT 425.310 499.610 425.690 499.620 ;
        RECT 424.880 499.310 425.690 499.610 ;
        RECT 425.310 499.300 425.690 499.310 ;
        RECT 425.335 499.295 425.665 499.300 ;
        RECT 425.310 496.890 425.690 496.900 ;
        RECT 426.025 496.890 426.355 496.905 ;
        RECT 425.310 496.590 426.355 496.890 ;
        RECT 425.310 496.580 425.690 496.590 ;
        RECT 426.025 496.575 426.355 496.590 ;
      LAYER via3 ;
        RECT 425.340 499.300 425.660 499.620 ;
        RECT 425.340 496.580 425.660 496.900 ;
      LAYER met4 ;
        RECT 425.335 499.295 425.665 499.625 ;
        RECT 425.350 496.905 425.650 499.295 ;
        RECT 425.335 496.575 425.665 496.905 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 426.720 498.820 427.040 499.080 ;
        RECT 426.810 498.680 426.950 498.820 ;
        RECT 426.810 498.540 427.180 498.680 ;
        RECT 427.040 498.400 427.180 498.540 ;
        RECT 426.950 498.140 427.270 498.400 ;
        RECT 282.970 438.500 283.290 438.560 ;
        RECT 427.410 438.500 427.730 438.560 ;
        RECT 282.970 438.360 427.730 438.500 ;
        RECT 282.970 438.300 283.290 438.360 ;
        RECT 427.410 438.300 427.730 438.360 ;
      LAYER via ;
        RECT 426.750 498.820 427.010 499.080 ;
        RECT 426.980 498.140 427.240 498.400 ;
        RECT 283.000 438.300 283.260 438.560 ;
        RECT 427.440 438.300 427.700 438.560 ;
      LAYER met2 ;
        RECT 426.770 500.000 427.050 504.000 ;
        RECT 426.810 499.110 426.950 500.000 ;
        RECT 426.750 498.790 427.010 499.110 ;
        RECT 426.980 498.110 427.240 498.430 ;
        RECT 427.040 483.070 427.180 498.110 ;
        RECT 427.040 482.930 427.640 483.070 ;
        RECT 427.500 438.590 427.640 482.930 ;
        RECT 283.000 438.270 283.260 438.590 ;
        RECT 427.440 438.270 427.700 438.590 ;
        RECT 283.060 82.870 283.200 438.270 ;
        RECT 283.060 82.730 286.880 82.870 ;
        RECT 286.740 2.400 286.880 82.730 ;
        RECT 286.530 -4.800 287.090 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.100 498.820 428.420 499.080 ;
        RECT 428.190 498.400 428.330 498.820 ;
        RECT 428.190 498.200 428.650 498.400 ;
        RECT 428.330 498.140 428.650 498.200 ;
        RECT 296.770 16.900 297.090 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 296.770 16.760 303.530 16.900 ;
        RECT 296.770 16.700 297.090 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 428.130 498.820 428.390 499.080 ;
        RECT 428.360 498.140 428.620 498.400 ;
        RECT 296.800 16.700 297.060 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 428.150 500.000 428.430 504.000 ;
        RECT 428.190 499.110 428.330 500.000 ;
        RECT 428.130 498.790 428.390 499.110 ;
        RECT 428.360 498.110 428.620 498.430 ;
        RECT 428.420 491.485 428.560 498.110 ;
        RECT 428.350 491.115 428.630 491.485 ;
        RECT 296.790 437.395 297.070 437.765 ;
        RECT 296.860 16.990 297.000 437.395 ;
        RECT 296.800 16.670 297.060 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 303.300 2.400 303.440 16.670 ;
        RECT 303.090 -4.800 303.650 2.400 ;
      LAYER via2 ;
        RECT 428.350 491.160 428.630 491.440 ;
        RECT 296.790 437.440 297.070 437.720 ;
      LAYER met3 ;
        RECT 428.325 491.450 428.655 491.465 ;
        RECT 428.990 491.450 429.370 491.460 ;
        RECT 428.325 491.150 429.370 491.450 ;
        RECT 428.325 491.135 428.655 491.150 ;
        RECT 428.990 491.140 429.370 491.150 ;
        RECT 296.765 437.730 297.095 437.745 ;
        RECT 428.990 437.730 429.370 437.740 ;
        RECT 296.765 437.430 429.370 437.730 ;
        RECT 296.765 437.415 297.095 437.430 ;
        RECT 428.990 437.420 429.370 437.430 ;
      LAYER via3 ;
        RECT 429.020 491.140 429.340 491.460 ;
        RECT 429.020 437.420 429.340 437.740 ;
      LAYER met4 ;
        RECT 429.015 491.135 429.345 491.465 ;
        RECT 429.030 437.745 429.330 491.135 ;
        RECT 429.015 437.415 429.345 437.745 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.480 499.160 429.800 499.420 ;
        RECT 429.570 498.340 429.710 499.160 ;
        RECT 430.170 498.340 430.490 498.400 ;
        RECT 429.570 498.200 430.490 498.340 ;
        RECT 430.170 498.140 430.490 498.200 ;
        RECT 319.770 32.540 320.090 32.600 ;
        RECT 430.630 32.540 430.950 32.600 ;
        RECT 319.770 32.400 430.950 32.540 ;
        RECT 319.770 32.340 320.090 32.400 ;
        RECT 430.630 32.340 430.950 32.400 ;
      LAYER via ;
        RECT 429.510 499.160 429.770 499.420 ;
        RECT 430.200 498.140 430.460 498.400 ;
        RECT 319.800 32.340 320.060 32.600 ;
        RECT 430.660 32.340 430.920 32.600 ;
      LAYER met2 ;
        RECT 429.530 500.000 429.810 504.000 ;
        RECT 429.570 499.450 429.710 500.000 ;
        RECT 429.510 499.130 429.770 499.450 ;
        RECT 430.200 498.110 430.460 498.430 ;
        RECT 430.260 472.840 430.400 498.110 ;
        RECT 430.260 472.700 430.860 472.840 ;
        RECT 430.720 32.630 430.860 472.700 ;
        RECT 319.800 32.310 320.060 32.630 ;
        RECT 430.660 32.310 430.920 32.630 ;
        RECT 319.860 2.400 320.000 32.310 ;
        RECT 319.650 -4.800 320.210 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 413.150 483.380 413.470 483.440 ;
        RECT 415.450 483.380 415.770 483.440 ;
        RECT 413.150 483.240 415.770 483.380 ;
        RECT 413.150 483.180 413.470 483.240 ;
        RECT 415.450 483.180 415.770 483.240 ;
        RECT 151.870 224.300 152.190 224.360 ;
        RECT 412.690 224.300 413.010 224.360 ;
        RECT 151.870 224.160 413.010 224.300 ;
        RECT 151.870 224.100 152.190 224.160 ;
        RECT 412.690 224.100 413.010 224.160 ;
      LAYER via ;
        RECT 413.180 483.180 413.440 483.440 ;
        RECT 415.480 483.180 415.740 483.440 ;
        RECT 151.900 224.100 152.160 224.360 ;
        RECT 412.720 224.100 412.980 224.360 ;
      LAYER met2 ;
        RECT 415.730 500.000 416.010 504.000 ;
        RECT 415.770 498.850 415.910 500.000 ;
        RECT 415.540 498.710 415.910 498.850 ;
        RECT 415.540 483.470 415.680 498.710 ;
        RECT 413.180 483.150 413.440 483.470 ;
        RECT 415.480 483.150 415.740 483.470 ;
        RECT 413.240 472.500 413.380 483.150 ;
        RECT 412.780 472.360 413.380 472.500 ;
        RECT 412.780 224.390 412.920 472.360 ;
        RECT 151.900 224.070 152.160 224.390 ;
        RECT 412.720 224.070 412.980 224.390 ;
        RECT 151.960 82.870 152.100 224.070 ;
        RECT 151.960 82.730 154.400 82.870 ;
        RECT 154.260 2.400 154.400 82.730 ;
        RECT 154.050 -4.800 154.610 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 431.320 499.500 431.640 499.760 ;
        RECT 431.410 499.080 431.550 499.500 ;
        RECT 431.410 498.880 431.870 499.080 ;
        RECT 431.550 498.820 431.870 498.880 ;
        RECT 341.850 33.220 342.170 33.280 ;
        RECT 430.170 33.220 430.490 33.280 ;
        RECT 341.850 33.080 430.490 33.220 ;
        RECT 341.850 33.020 342.170 33.080 ;
        RECT 430.170 33.020 430.490 33.080 ;
      LAYER via ;
        RECT 431.350 499.500 431.610 499.760 ;
        RECT 431.580 498.820 431.840 499.080 ;
        RECT 341.880 33.020 342.140 33.280 ;
        RECT 430.200 33.020 430.460 33.280 ;
      LAYER met2 ;
        RECT 431.370 500.000 431.650 504.000 ;
        RECT 431.410 499.790 431.550 500.000 ;
        RECT 431.350 499.470 431.610 499.790 ;
        RECT 431.580 498.965 431.840 499.110 ;
        RECT 431.570 498.595 431.850 498.965 ;
        RECT 429.730 497.915 430.010 498.285 ;
        RECT 429.800 472.500 429.940 497.915 ;
        RECT 429.800 472.360 430.400 472.500 ;
        RECT 430.260 33.310 430.400 472.360 ;
        RECT 341.880 32.990 342.140 33.310 ;
        RECT 430.200 32.990 430.460 33.310 ;
        RECT 341.940 2.400 342.080 32.990 ;
        RECT 341.730 -4.800 342.290 2.400 ;
      LAYER via2 ;
        RECT 431.570 498.640 431.850 498.920 ;
        RECT 429.730 497.960 430.010 498.240 ;
      LAYER met3 ;
        RECT 431.545 498.930 431.875 498.945 ;
        RECT 430.870 498.630 431.875 498.930 ;
        RECT 429.705 498.250 430.035 498.265 ;
        RECT 430.870 498.250 431.170 498.630 ;
        RECT 431.545 498.615 431.875 498.630 ;
        RECT 429.705 497.950 431.170 498.250 ;
        RECT 429.705 497.935 430.035 497.950 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.930 499.160 433.250 499.420 ;
        RECT 433.020 498.740 433.160 499.160 ;
        RECT 432.930 498.480 433.250 498.740 ;
        RECT 413.610 491.540 413.930 491.600 ;
        RECT 432.930 491.540 433.250 491.600 ;
        RECT 413.610 491.400 433.250 491.540 ;
        RECT 413.610 491.340 413.930 491.400 ;
        RECT 432.930 491.340 433.250 491.400 ;
        RECT 351.970 224.980 352.290 225.040 ;
        RECT 413.150 224.980 413.470 225.040 ;
        RECT 351.970 224.840 413.470 224.980 ;
        RECT 351.970 224.780 352.290 224.840 ;
        RECT 413.150 224.780 413.470 224.840 ;
        RECT 351.970 16.900 352.290 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 351.970 16.760 358.730 16.900 ;
        RECT 351.970 16.700 352.290 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 432.960 499.160 433.220 499.420 ;
        RECT 432.960 498.480 433.220 498.740 ;
        RECT 413.640 491.340 413.900 491.600 ;
        RECT 432.960 491.340 433.220 491.600 ;
        RECT 352.000 224.780 352.260 225.040 ;
        RECT 413.180 224.780 413.440 225.040 ;
        RECT 352.000 16.700 352.260 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 432.750 500.000 433.030 504.000 ;
        RECT 432.790 499.530 432.930 500.000 ;
        RECT 432.790 499.450 433.160 499.530 ;
        RECT 432.790 499.390 433.220 499.450 ;
        RECT 432.960 499.130 433.220 499.390 ;
        RECT 432.960 498.450 433.220 498.770 ;
        RECT 433.020 491.630 433.160 498.450 ;
        RECT 413.640 491.310 413.900 491.630 ;
        RECT 432.960 491.310 433.220 491.630 ;
        RECT 413.700 448.570 413.840 491.310 ;
        RECT 413.240 448.430 413.840 448.570 ;
        RECT 413.240 225.070 413.380 448.430 ;
        RECT 352.000 224.750 352.260 225.070 ;
        RECT 413.180 224.750 413.440 225.070 ;
        RECT 352.060 16.990 352.200 224.750 ;
        RECT 352.000 16.670 352.260 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 358.500 2.400 358.640 16.670 ;
        RECT 358.290 -4.800 358.850 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.250 472.160 429.570 472.220 ;
        RECT 434.310 472.160 434.630 472.220 ;
        RECT 429.250 472.020 434.630 472.160 ;
        RECT 429.250 471.960 429.570 472.020 ;
        RECT 434.310 471.960 434.630 472.020 ;
        RECT 374.970 26.760 375.290 26.820 ;
        RECT 429.250 26.760 429.570 26.820 ;
        RECT 374.970 26.620 429.570 26.760 ;
        RECT 374.970 26.560 375.290 26.620 ;
        RECT 429.250 26.560 429.570 26.620 ;
      LAYER via ;
        RECT 429.280 471.960 429.540 472.220 ;
        RECT 434.340 471.960 434.600 472.220 ;
        RECT 375.000 26.560 375.260 26.820 ;
        RECT 429.280 26.560 429.540 26.820 ;
      LAYER met2 ;
        RECT 434.130 500.000 434.410 504.000 ;
        RECT 434.170 499.645 434.310 500.000 ;
        RECT 434.100 499.275 434.380 499.645 ;
        RECT 434.330 497.915 434.610 498.285 ;
        RECT 434.400 472.250 434.540 497.915 ;
        RECT 429.280 471.930 429.540 472.250 ;
        RECT 434.340 471.930 434.600 472.250 ;
        RECT 429.340 26.850 429.480 471.930 ;
        RECT 375.000 26.530 375.260 26.850 ;
        RECT 429.280 26.530 429.540 26.850 ;
        RECT 375.060 2.400 375.200 26.530 ;
        RECT 374.850 -4.800 375.410 2.400 ;
      LAYER via2 ;
        RECT 434.100 499.320 434.380 499.600 ;
        RECT 434.330 497.960 434.610 498.240 ;
      LAYER met3 ;
        RECT 434.075 499.610 434.405 499.625 ;
        RECT 432.710 499.310 434.405 499.610 ;
        RECT 432.710 498.250 433.010 499.310 ;
        RECT 434.075 499.295 434.405 499.310 ;
        RECT 434.305 498.250 434.635 498.265 ;
        RECT 432.710 497.950 434.635 498.250 ;
        RECT 434.305 497.935 434.635 497.950 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.690 473.320 436.010 473.580 ;
        RECT 435.780 473.180 435.920 473.320 ;
        RECT 435.780 473.040 440.980 473.180 ;
        RECT 440.290 471.820 440.610 471.880 ;
        RECT 440.840 471.820 440.980 473.040 ;
        RECT 440.290 471.680 440.980 471.820 ;
        RECT 440.290 471.620 440.610 471.680 ;
        RECT 386.470 438.840 386.790 438.900 ;
        RECT 440.290 438.840 440.610 438.900 ;
        RECT 386.470 438.700 440.610 438.840 ;
        RECT 386.470 438.640 386.790 438.700 ;
        RECT 440.290 438.640 440.610 438.700 ;
      LAYER via ;
        RECT 435.720 473.320 435.980 473.580 ;
        RECT 440.320 471.620 440.580 471.880 ;
        RECT 386.500 438.640 386.760 438.900 ;
        RECT 440.320 438.640 440.580 438.900 ;
      LAYER met2 ;
        RECT 435.510 500.000 435.790 504.000 ;
        RECT 435.550 499.020 435.690 500.000 ;
        RECT 435.320 498.880 435.690 499.020 ;
        RECT 435.320 497.320 435.460 498.880 ;
        RECT 435.320 497.180 435.920 497.320 ;
        RECT 435.780 473.610 435.920 497.180 ;
        RECT 435.720 473.290 435.980 473.610 ;
        RECT 440.320 471.590 440.580 471.910 ;
        RECT 440.380 438.930 440.520 471.590 ;
        RECT 386.500 438.610 386.760 438.930 ;
        RECT 440.320 438.610 440.580 438.930 ;
        RECT 386.560 82.870 386.700 438.610 ;
        RECT 386.560 82.730 391.760 82.870 ;
        RECT 391.620 2.400 391.760 82.730 ;
        RECT 391.410 -4.800 391.970 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 409.010 485.420 409.330 485.480 ;
        RECT 438.910 485.420 439.230 485.480 ;
        RECT 409.010 485.280 439.230 485.420 ;
        RECT 409.010 485.220 409.330 485.280 ;
        RECT 438.910 485.220 439.230 485.280 ;
      LAYER via ;
        RECT 409.040 485.220 409.300 485.480 ;
        RECT 438.940 485.220 439.200 485.480 ;
      LAYER met2 ;
        RECT 436.890 500.000 437.170 504.000 ;
        RECT 436.930 498.850 437.070 500.000 ;
        RECT 436.930 498.710 437.300 498.850 ;
        RECT 437.160 498.285 437.300 498.710 ;
        RECT 437.090 497.915 437.370 498.285 ;
        RECT 438.930 497.235 439.210 497.605 ;
        RECT 439.000 485.510 439.140 497.235 ;
        RECT 409.040 485.190 409.300 485.510 ;
        RECT 438.940 485.190 439.200 485.510 ;
        RECT 407.970 1.770 408.530 2.400 ;
        RECT 409.100 1.770 409.240 485.190 ;
        RECT 407.970 1.630 409.240 1.770 ;
        RECT 407.970 -4.800 408.530 1.630 ;
      LAYER via2 ;
        RECT 437.090 497.960 437.370 498.240 ;
        RECT 438.930 497.280 439.210 497.560 ;
      LAYER met3 ;
        RECT 437.065 498.250 437.395 498.265 ;
        RECT 437.065 497.950 439.220 498.250 ;
        RECT 437.065 497.935 437.395 497.950 ;
        RECT 438.920 497.585 439.220 497.950 ;
        RECT 438.905 497.255 439.235 497.585 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.730 100.200 424.050 100.260 ;
        RECT 438.910 100.200 439.230 100.260 ;
        RECT 423.730 100.060 439.230 100.200 ;
        RECT 423.730 100.000 424.050 100.060 ;
        RECT 438.910 100.000 439.230 100.060 ;
      LAYER via ;
        RECT 423.760 100.000 424.020 100.260 ;
        RECT 438.940 100.000 439.200 100.260 ;
      LAYER met2 ;
        RECT 438.270 500.000 438.550 504.000 ;
        RECT 438.310 498.340 438.450 500.000 ;
        RECT 438.310 498.200 438.680 498.340 ;
        RECT 438.540 476.170 438.680 498.200 ;
        RECT 438.540 476.030 439.140 476.170 ;
        RECT 439.000 100.290 439.140 476.030 ;
        RECT 423.760 99.970 424.020 100.290 ;
        RECT 438.940 99.970 439.200 100.290 ;
        RECT 423.820 17.410 423.960 99.970 ;
        RECT 423.820 17.270 424.880 17.410 ;
        RECT 424.740 2.400 424.880 17.270 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.650 500.000 439.930 504.000 ;
        RECT 439.690 499.020 439.830 500.000 ;
        RECT 439.690 498.965 440.520 499.020 ;
        RECT 439.690 498.880 440.590 498.965 ;
        RECT 440.310 498.595 440.590 498.880 ;
        RECT 440.770 497.235 441.050 497.605 ;
        RECT 440.840 82.870 440.980 497.235 ;
        RECT 440.840 82.730 441.440 82.870 ;
        RECT 441.300 2.400 441.440 82.730 ;
        RECT 441.090 -4.800 441.650 2.400 ;
      LAYER via2 ;
        RECT 440.310 498.640 440.590 498.920 ;
        RECT 440.770 497.280 441.050 497.560 ;
      LAYER met3 ;
        RECT 440.285 498.930 440.615 498.945 ;
        RECT 440.285 498.630 441.290 498.930 ;
        RECT 440.285 498.615 440.615 498.630 ;
        RECT 440.990 497.585 441.290 498.630 ;
        RECT 440.745 497.270 441.290 497.585 ;
        RECT 440.745 497.255 441.075 497.270 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 440.750 497.800 441.070 498.060 ;
        RECT 440.840 496.980 440.980 497.800 ;
        RECT 446.730 496.980 447.050 497.040 ;
        RECT 440.840 496.840 447.050 496.980 ;
        RECT 446.730 496.780 447.050 496.840 ;
        RECT 446.730 17.580 447.050 17.640 ;
        RECT 457.770 17.580 458.090 17.640 ;
        RECT 446.730 17.440 458.090 17.580 ;
        RECT 446.730 17.380 447.050 17.440 ;
        RECT 457.770 17.380 458.090 17.440 ;
      LAYER via ;
        RECT 440.780 497.800 441.040 498.060 ;
        RECT 446.760 496.780 447.020 497.040 ;
        RECT 446.760 17.380 447.020 17.640 ;
        RECT 457.800 17.380 458.060 17.640 ;
      LAYER met2 ;
        RECT 441.030 500.000 441.310 504.000 ;
        RECT 441.070 498.680 441.210 500.000 ;
        RECT 440.840 498.540 441.210 498.680 ;
        RECT 440.840 498.090 440.980 498.540 ;
        RECT 440.780 497.770 441.040 498.090 ;
        RECT 446.760 496.750 447.020 497.070 ;
        RECT 446.820 17.670 446.960 496.750 ;
        RECT 446.760 17.350 447.020 17.670 ;
        RECT 457.800 17.350 458.060 17.670 ;
        RECT 457.860 2.400 458.000 17.350 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.360 499.500 442.680 499.760 ;
        RECT 442.450 499.020 442.590 499.500 ;
        RECT 442.450 498.880 443.050 499.020 ;
        RECT 442.130 497.320 442.450 497.380 ;
        RECT 442.910 497.320 443.050 498.880 ;
        RECT 442.130 497.180 443.050 497.320 ;
        RECT 442.130 497.120 442.450 497.180 ;
        RECT 443.510 21.660 443.830 21.720 ;
        RECT 474.330 21.660 474.650 21.720 ;
        RECT 443.510 21.520 474.650 21.660 ;
        RECT 443.510 21.460 443.830 21.520 ;
        RECT 474.330 21.460 474.650 21.520 ;
      LAYER via ;
        RECT 442.390 499.500 442.650 499.760 ;
        RECT 442.160 497.120 442.420 497.380 ;
        RECT 443.540 21.460 443.800 21.720 ;
        RECT 474.360 21.460 474.620 21.720 ;
      LAYER met2 ;
        RECT 442.410 500.000 442.690 504.000 ;
        RECT 442.450 499.790 442.590 500.000 ;
        RECT 442.390 499.470 442.650 499.790 ;
        RECT 442.160 497.090 442.420 497.410 ;
        RECT 442.220 488.650 442.360 497.090 ;
        RECT 442.220 488.510 442.820 488.650 ;
        RECT 442.680 472.500 442.820 488.510 ;
        RECT 442.680 472.360 443.740 472.500 ;
        RECT 443.600 21.750 443.740 472.360 ;
        RECT 443.540 21.430 443.800 21.750 ;
        RECT 474.360 21.430 474.620 21.750 ;
        RECT 474.420 2.400 474.560 21.430 ;
        RECT 474.210 -4.800 474.770 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.740 499.360 444.060 499.420 ;
        RECT 443.370 499.220 444.060 499.360 ;
        RECT 443.370 497.380 443.510 499.220 ;
        RECT 443.740 499.160 444.060 499.220 ;
        RECT 443.370 497.180 443.830 497.380 ;
        RECT 443.510 497.120 443.830 497.180 ;
        RECT 443.510 473.860 443.830 473.920 ;
        RECT 445.350 473.860 445.670 473.920 ;
        RECT 443.510 473.720 445.670 473.860 ;
        RECT 443.510 473.660 443.830 473.720 ;
        RECT 445.350 473.660 445.670 473.720 ;
        RECT 445.350 99.860 445.670 99.920 ;
        RECT 490.430 99.860 490.750 99.920 ;
        RECT 445.350 99.720 490.750 99.860 ;
        RECT 445.350 99.660 445.670 99.720 ;
        RECT 490.430 99.660 490.750 99.720 ;
      LAYER via ;
        RECT 443.770 499.160 444.030 499.420 ;
        RECT 443.540 497.120 443.800 497.380 ;
        RECT 443.540 473.660 443.800 473.920 ;
        RECT 445.380 473.660 445.640 473.920 ;
        RECT 445.380 99.660 445.640 99.920 ;
        RECT 490.460 99.660 490.720 99.920 ;
      LAYER met2 ;
        RECT 443.790 500.000 444.070 504.000 ;
        RECT 443.830 499.450 443.970 500.000 ;
        RECT 443.770 499.130 444.030 499.450 ;
        RECT 443.540 497.090 443.800 497.410 ;
        RECT 443.600 473.950 443.740 497.090 ;
        RECT 443.540 473.630 443.800 473.950 ;
        RECT 445.380 473.630 445.640 473.950 ;
        RECT 445.440 99.950 445.580 473.630 ;
        RECT 445.380 99.630 445.640 99.950 ;
        RECT 490.460 99.630 490.720 99.950 ;
        RECT 490.520 82.870 490.660 99.630 ;
        RECT 490.520 82.730 491.120 82.870 ;
        RECT 490.980 2.400 491.120 82.730 ;
        RECT 490.770 -4.800 491.330 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 417.520 499.700 417.840 499.760 ;
        RECT 413.470 499.560 417.840 499.700 ;
        RECT 398.890 498.680 399.210 498.740 ;
        RECT 413.470 498.680 413.610 499.560 ;
        RECT 417.520 499.500 417.840 499.560 ;
        RECT 398.890 498.540 413.610 498.680 ;
        RECT 398.890 498.480 399.210 498.540 ;
        RECT 265.490 487.460 265.810 487.520 ;
        RECT 398.890 487.460 399.210 487.520 ;
        RECT 265.490 487.320 399.210 487.460 ;
        RECT 265.490 487.260 265.810 487.320 ;
        RECT 398.890 487.260 399.210 487.320 ;
        RECT 176.250 18.940 176.570 19.000 ;
        RECT 265.490 18.940 265.810 19.000 ;
        RECT 176.250 18.800 265.810 18.940 ;
        RECT 176.250 18.740 176.570 18.800 ;
        RECT 265.490 18.740 265.810 18.800 ;
      LAYER via ;
        RECT 398.920 498.480 399.180 498.740 ;
        RECT 417.550 499.500 417.810 499.760 ;
        RECT 265.520 487.260 265.780 487.520 ;
        RECT 398.920 487.260 399.180 487.520 ;
        RECT 176.280 18.740 176.540 19.000 ;
        RECT 265.520 18.740 265.780 19.000 ;
      LAYER met2 ;
        RECT 417.570 500.000 417.850 504.000 ;
        RECT 417.610 499.790 417.750 500.000 ;
        RECT 417.550 499.470 417.810 499.790 ;
        RECT 398.920 498.450 399.180 498.770 ;
        RECT 398.980 487.550 399.120 498.450 ;
        RECT 265.520 487.230 265.780 487.550 ;
        RECT 398.920 487.230 399.180 487.550 ;
        RECT 265.580 19.030 265.720 487.230 ;
        RECT 176.280 18.710 176.540 19.030 ;
        RECT 265.520 18.710 265.780 19.030 ;
        RECT 176.340 2.400 176.480 18.710 ;
        RECT 176.130 -4.800 176.690 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 231.440 446.130 231.500 ;
        RECT 500.090 231.440 500.410 231.500 ;
        RECT 445.810 231.300 500.410 231.440 ;
        RECT 445.810 231.240 446.130 231.300 ;
        RECT 500.090 231.240 500.410 231.300 ;
        RECT 500.090 16.900 500.410 16.960 ;
        RECT 507.450 16.900 507.770 16.960 ;
        RECT 500.090 16.760 507.770 16.900 ;
        RECT 500.090 16.700 500.410 16.760 ;
        RECT 507.450 16.700 507.770 16.760 ;
      LAYER via ;
        RECT 445.840 231.240 446.100 231.500 ;
        RECT 500.120 231.240 500.380 231.500 ;
        RECT 500.120 16.700 500.380 16.960 ;
        RECT 507.480 16.700 507.740 16.960 ;
      LAYER met2 ;
        RECT 445.170 500.000 445.450 504.000 ;
        RECT 445.210 498.850 445.350 500.000 ;
        RECT 445.210 498.710 445.580 498.850 ;
        RECT 445.440 498.170 445.580 498.710 ;
        RECT 445.440 498.030 446.040 498.170 ;
        RECT 445.900 231.530 446.040 498.030 ;
        RECT 445.840 231.210 446.100 231.530 ;
        RECT 500.120 231.210 500.380 231.530 ;
        RECT 500.180 16.990 500.320 231.210 ;
        RECT 500.120 16.670 500.380 16.990 ;
        RECT 507.480 16.670 507.740 16.990 ;
        RECT 507.540 2.400 507.680 16.670 ;
        RECT 507.330 -4.800 507.890 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.500 499.500 446.820 499.760 ;
        RECT 446.590 498.000 446.730 499.500 ;
        RECT 446.590 497.860 449.720 498.000 ;
        RECT 449.580 497.720 449.720 497.860 ;
        RECT 449.490 497.460 449.810 497.720 ;
        RECT 472.490 19.620 472.810 19.680 ;
        RECT 524.010 19.620 524.330 19.680 ;
        RECT 472.490 19.480 524.330 19.620 ;
        RECT 472.490 19.420 472.810 19.480 ;
        RECT 524.010 19.420 524.330 19.480 ;
      LAYER via ;
        RECT 446.530 499.500 446.790 499.760 ;
        RECT 449.520 497.460 449.780 497.720 ;
        RECT 472.520 19.420 472.780 19.680 ;
        RECT 524.040 19.420 524.300 19.680 ;
      LAYER met2 ;
        RECT 446.550 500.000 446.830 504.000 ;
        RECT 446.590 499.790 446.730 500.000 ;
        RECT 446.530 499.470 446.790 499.790 ;
        RECT 449.520 497.430 449.780 497.750 ;
        RECT 449.580 492.165 449.720 497.430 ;
        RECT 449.510 491.795 449.790 492.165 ;
        RECT 472.510 440.795 472.790 441.165 ;
        RECT 472.580 19.710 472.720 440.795 ;
        RECT 472.520 19.390 472.780 19.710 ;
        RECT 524.040 19.390 524.300 19.710 ;
        RECT 524.100 2.400 524.240 19.390 ;
        RECT 523.890 -4.800 524.450 2.400 ;
      LAYER via2 ;
        RECT 449.510 491.840 449.790 492.120 ;
        RECT 472.510 440.840 472.790 441.120 ;
      LAYER met3 ;
        RECT 446.470 492.130 446.850 492.140 ;
        RECT 449.485 492.130 449.815 492.145 ;
        RECT 446.470 491.830 449.815 492.130 ;
        RECT 446.470 491.820 446.850 491.830 ;
        RECT 449.485 491.815 449.815 491.830 ;
        RECT 446.470 441.130 446.850 441.140 ;
        RECT 472.485 441.130 472.815 441.145 ;
        RECT 446.470 440.830 472.815 441.130 ;
        RECT 446.470 440.820 446.850 440.830 ;
        RECT 472.485 440.815 472.815 440.830 ;
      LAYER via3 ;
        RECT 446.500 491.820 446.820 492.140 ;
        RECT 446.500 440.820 446.820 441.140 ;
      LAYER met4 ;
        RECT 446.495 491.815 446.825 492.145 ;
        RECT 446.510 441.145 446.810 491.815 ;
        RECT 446.495 440.815 446.825 441.145 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 447.880 499.500 448.200 499.760 ;
        RECT 447.970 498.400 448.110 499.500 ;
        RECT 447.650 498.200 448.110 498.400 ;
        RECT 447.650 498.140 447.970 498.200 ;
        RECT 447.650 485.760 447.970 485.820 ;
        RECT 452.250 485.760 452.570 485.820 ;
        RECT 447.650 485.620 452.570 485.760 ;
        RECT 447.650 485.560 447.970 485.620 ;
        RECT 452.250 485.560 452.570 485.620 ;
        RECT 452.250 25.740 452.570 25.800 ;
        RECT 452.250 25.600 479.160 25.740 ;
        RECT 452.250 25.540 452.570 25.600 ;
        RECT 479.020 25.400 479.160 25.600 ;
        RECT 479.020 25.260 493.420 25.400 ;
        RECT 493.280 25.060 493.420 25.260 ;
        RECT 540.570 25.060 540.890 25.120 ;
        RECT 493.280 24.920 540.890 25.060 ;
        RECT 540.570 24.860 540.890 24.920 ;
      LAYER via ;
        RECT 447.910 499.500 448.170 499.760 ;
        RECT 447.680 498.140 447.940 498.400 ;
        RECT 447.680 485.560 447.940 485.820 ;
        RECT 452.280 485.560 452.540 485.820 ;
        RECT 452.280 25.540 452.540 25.800 ;
        RECT 540.600 24.860 540.860 25.120 ;
      LAYER met2 ;
        RECT 447.930 500.000 448.210 504.000 ;
        RECT 447.970 499.790 448.110 500.000 ;
        RECT 447.910 499.470 448.170 499.790 ;
        RECT 447.680 498.110 447.940 498.430 ;
        RECT 447.740 485.850 447.880 498.110 ;
        RECT 447.680 485.530 447.940 485.850 ;
        RECT 452.280 485.530 452.540 485.850 ;
        RECT 452.340 25.830 452.480 485.530 ;
        RECT 452.280 25.510 452.540 25.830 ;
        RECT 540.600 24.830 540.860 25.150 ;
        RECT 540.660 2.400 540.800 24.830 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 472.160 449.350 472.220 ;
        RECT 451.330 472.160 451.650 472.220 ;
        RECT 449.030 472.020 451.650 472.160 ;
        RECT 449.030 471.960 449.350 472.020 ;
        RECT 451.330 471.960 451.650 472.020 ;
        RECT 451.330 107.000 451.650 107.060 ;
        RECT 552.990 107.000 553.310 107.060 ;
        RECT 451.330 106.860 553.310 107.000 ;
        RECT 451.330 106.800 451.650 106.860 ;
        RECT 552.990 106.800 553.310 106.860 ;
      LAYER via ;
        RECT 449.060 471.960 449.320 472.220 ;
        RECT 451.360 471.960 451.620 472.220 ;
        RECT 451.360 106.800 451.620 107.060 ;
        RECT 553.020 106.800 553.280 107.060 ;
      LAYER met2 ;
        RECT 449.310 500.000 449.590 504.000 ;
        RECT 449.350 499.815 449.490 500.000 ;
        RECT 449.280 499.445 449.560 499.815 ;
        RECT 449.050 497.915 449.330 498.285 ;
        RECT 449.120 472.250 449.260 497.915 ;
        RECT 449.060 471.930 449.320 472.250 ;
        RECT 451.360 471.930 451.620 472.250 ;
        RECT 451.420 107.090 451.560 471.930 ;
        RECT 451.360 106.770 451.620 107.090 ;
        RECT 553.020 106.770 553.280 107.090 ;
        RECT 553.080 82.870 553.220 106.770 ;
        RECT 553.080 82.730 557.360 82.870 ;
        RECT 557.220 2.400 557.360 82.730 ;
        RECT 557.010 -4.800 557.570 2.400 ;
      LAYER via2 ;
        RECT 449.280 499.490 449.560 499.770 ;
        RECT 449.050 497.960 449.330 498.240 ;
      LAYER met3 ;
        RECT 449.255 499.465 449.585 499.795 ;
        RECT 449.270 498.265 449.570 499.465 ;
        RECT 449.025 497.950 449.570 498.265 ;
        RECT 449.025 497.935 449.355 497.950 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 450.410 490.520 450.730 490.580 ;
        RECT 458.690 490.520 459.010 490.580 ;
        RECT 450.410 490.380 459.010 490.520 ;
        RECT 450.410 490.320 450.730 490.380 ;
        RECT 458.690 490.320 459.010 490.380 ;
        RECT 458.690 31.520 459.010 31.580 ;
        RECT 573.690 31.520 574.010 31.580 ;
        RECT 458.690 31.380 574.010 31.520 ;
        RECT 458.690 31.320 459.010 31.380 ;
        RECT 573.690 31.320 574.010 31.380 ;
      LAYER via ;
        RECT 450.440 490.320 450.700 490.580 ;
        RECT 458.720 490.320 458.980 490.580 ;
        RECT 458.720 31.320 458.980 31.580 ;
        RECT 573.720 31.320 573.980 31.580 ;
      LAYER met2 ;
        RECT 450.690 500.000 450.970 504.000 ;
        RECT 450.730 498.340 450.870 500.000 ;
        RECT 450.500 498.200 450.870 498.340 ;
        RECT 450.500 490.610 450.640 498.200 ;
        RECT 450.440 490.290 450.700 490.610 ;
        RECT 458.720 490.290 458.980 490.610 ;
        RECT 458.780 31.610 458.920 490.290 ;
        RECT 458.720 31.290 458.980 31.610 ;
        RECT 573.720 31.290 573.980 31.610 ;
        RECT 573.780 2.400 573.920 31.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 452.020 499.500 452.340 499.760 ;
        RECT 452.110 499.360 452.250 499.500 ;
        RECT 452.110 499.220 452.940 499.360 ;
        RECT 452.800 498.400 452.940 499.220 ;
        RECT 452.710 498.140 453.030 498.400 ;
        RECT 449.030 471.480 449.350 471.540 ;
        RECT 452.710 471.480 453.030 471.540 ;
        RECT 449.030 471.340 453.030 471.480 ;
        RECT 449.030 471.280 449.350 471.340 ;
        RECT 452.710 471.280 453.030 471.340 ;
        RECT 590.250 17.240 590.570 17.300 ;
        RECT 469.130 17.100 590.570 17.240 ;
        RECT 449.030 16.560 449.350 16.620 ;
        RECT 469.130 16.560 469.270 17.100 ;
        RECT 590.250 17.040 590.570 17.100 ;
        RECT 449.030 16.420 469.270 16.560 ;
        RECT 449.030 16.360 449.350 16.420 ;
      LAYER via ;
        RECT 452.050 499.500 452.310 499.760 ;
        RECT 452.740 498.140 453.000 498.400 ;
        RECT 449.060 471.280 449.320 471.540 ;
        RECT 452.740 471.280 453.000 471.540 ;
        RECT 449.060 16.360 449.320 16.620 ;
        RECT 590.280 17.040 590.540 17.300 ;
      LAYER met2 ;
        RECT 452.070 500.000 452.350 504.000 ;
        RECT 452.110 499.790 452.250 500.000 ;
        RECT 452.050 499.470 452.310 499.790 ;
        RECT 452.740 498.110 453.000 498.430 ;
        RECT 452.800 471.570 452.940 498.110 ;
        RECT 449.060 471.250 449.320 471.570 ;
        RECT 452.740 471.250 453.000 471.570 ;
        RECT 449.120 16.650 449.260 471.250 ;
        RECT 590.280 17.010 590.540 17.330 ;
        RECT 449.060 16.330 449.320 16.650 ;
        RECT 590.340 2.400 590.480 17.010 ;
        RECT 590.130 -4.800 590.690 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.790 458.900 452.110 458.960 ;
        RECT 601.290 458.900 601.610 458.960 ;
        RECT 451.790 458.760 601.610 458.900 ;
        RECT 451.790 458.700 452.110 458.760 ;
        RECT 601.290 458.700 601.610 458.760 ;
      LAYER via ;
        RECT 451.820 458.700 452.080 458.960 ;
        RECT 601.320 458.700 601.580 458.960 ;
      LAYER met2 ;
        RECT 453.450 500.000 453.730 504.000 ;
        RECT 453.490 499.645 453.630 500.000 ;
        RECT 453.420 499.275 453.700 499.645 ;
        RECT 451.810 497.915 452.090 498.285 ;
        RECT 451.880 458.990 452.020 497.915 ;
        RECT 451.820 458.670 452.080 458.990 ;
        RECT 601.320 458.670 601.580 458.990 ;
        RECT 601.380 82.870 601.520 458.670 ;
        RECT 601.380 82.730 606.120 82.870 ;
        RECT 605.980 17.410 606.120 82.730 ;
        RECT 605.980 17.270 607.040 17.410 ;
        RECT 606.900 2.400 607.040 17.270 ;
        RECT 606.690 -4.800 607.250 2.400 ;
      LAYER via2 ;
        RECT 453.420 499.320 453.700 499.600 ;
        RECT 451.810 497.960 452.090 498.240 ;
      LAYER met3 ;
        RECT 453.395 499.610 453.725 499.625 ;
        RECT 452.030 499.310 453.725 499.610 ;
        RECT 452.030 498.265 452.330 499.310 ;
        RECT 453.395 499.295 453.725 499.310 ;
        RECT 451.785 497.950 452.330 498.265 ;
        RECT 451.785 497.935 452.115 497.950 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.830 500.000 455.110 504.000 ;
        RECT 454.870 499.815 455.010 500.000 ;
        RECT 454.800 499.445 455.080 499.815 ;
        RECT 623.390 16.475 623.670 16.845 ;
        RECT 623.460 2.400 623.600 16.475 ;
        RECT 623.250 -4.800 623.810 2.400 ;
      LAYER via2 ;
        RECT 454.800 499.490 455.080 499.770 ;
        RECT 623.390 16.520 623.670 16.800 ;
      LAYER met3 ;
        RECT 454.775 499.620 455.105 499.795 ;
        RECT 454.750 499.610 455.130 499.620 ;
        RECT 454.750 499.310 455.390 499.610 ;
        RECT 454.750 499.300 455.130 499.310 ;
        RECT 454.750 16.810 455.130 16.820 ;
        RECT 623.365 16.810 623.695 16.825 ;
        RECT 454.750 16.510 623.695 16.810 ;
        RECT 454.750 16.500 455.130 16.510 ;
        RECT 623.365 16.495 623.695 16.510 ;
      LAYER via3 ;
        RECT 454.780 499.300 455.100 499.620 ;
        RECT 454.780 16.500 455.100 16.820 ;
      LAYER met4 ;
        RECT 454.775 499.295 455.105 499.625 ;
        RECT 454.790 16.825 455.090 499.295 ;
        RECT 454.775 16.495 455.105 16.825 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.160 499.500 456.480 499.760 ;
        RECT 456.250 498.680 456.390 499.500 ;
        RECT 455.560 498.540 456.390 498.680 ;
        RECT 455.560 498.000 455.700 498.540 ;
        RECT 456.390 498.000 456.710 498.060 ;
        RECT 455.560 497.860 456.710 498.000 ;
        RECT 456.390 497.800 456.710 497.860 ;
        RECT 634.870 475.220 635.190 475.280 ;
        RECT 593.330 475.080 635.190 475.220 ;
        RECT 456.390 474.880 456.710 474.940 ;
        RECT 593.330 474.880 593.470 475.080 ;
        RECT 634.870 475.020 635.190 475.080 ;
        RECT 456.390 474.740 593.470 474.880 ;
        RECT 456.390 474.680 456.710 474.740 ;
      LAYER via ;
        RECT 456.190 499.500 456.450 499.760 ;
        RECT 456.420 497.800 456.680 498.060 ;
        RECT 456.420 474.680 456.680 474.940 ;
        RECT 634.900 475.020 635.160 475.280 ;
      LAYER met2 ;
        RECT 456.210 500.000 456.490 504.000 ;
        RECT 456.250 499.790 456.390 500.000 ;
        RECT 456.190 499.470 456.450 499.790 ;
        RECT 456.420 497.770 456.680 498.090 ;
        RECT 456.480 474.970 456.620 497.770 ;
        RECT 634.900 474.990 635.160 475.310 ;
        RECT 456.420 474.650 456.680 474.970 ;
        RECT 634.960 82.870 635.100 474.990 ;
        RECT 634.960 82.730 637.400 82.870 ;
        RECT 637.260 17.410 637.400 82.730 ;
        RECT 637.260 17.270 640.160 17.410 ;
        RECT 640.020 2.400 640.160 17.270 ;
        RECT 639.810 -4.800 640.370 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.540 499.160 457.860 499.420 ;
        RECT 457.630 497.660 457.770 499.160 ;
        RECT 461.450 497.660 461.770 497.720 ;
        RECT 457.630 497.520 461.770 497.660 ;
        RECT 461.450 497.460 461.770 497.520 ;
        RECT 461.910 489.500 462.230 489.560 ;
        RECT 461.910 489.360 496.870 489.500 ;
        RECT 461.910 489.300 462.230 489.360 ;
        RECT 496.730 489.160 496.870 489.360 ;
        RECT 655.570 489.160 655.890 489.220 ;
        RECT 496.730 489.020 655.890 489.160 ;
        RECT 655.570 488.960 655.890 489.020 ;
      LAYER via ;
        RECT 457.570 499.160 457.830 499.420 ;
        RECT 461.480 497.460 461.740 497.720 ;
        RECT 461.940 489.300 462.200 489.560 ;
        RECT 655.600 488.960 655.860 489.220 ;
      LAYER met2 ;
        RECT 457.590 500.000 457.870 504.000 ;
        RECT 457.630 499.450 457.770 500.000 ;
        RECT 457.570 499.130 457.830 499.450 ;
        RECT 461.480 497.660 461.740 497.750 ;
        RECT 461.480 497.520 462.140 497.660 ;
        RECT 461.480 497.430 461.740 497.520 ;
        RECT 462.000 489.590 462.140 497.520 ;
        RECT 461.940 489.270 462.200 489.590 ;
        RECT 655.600 488.930 655.860 489.250 ;
        RECT 655.660 17.410 655.800 488.930 ;
        RECT 655.660 17.270 656.720 17.410 ;
        RECT 656.580 2.400 656.720 17.270 ;
        RECT 656.370 -4.800 656.930 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 193.270 107.000 193.590 107.060 ;
        RECT 418.210 107.000 418.530 107.060 ;
        RECT 193.270 106.860 418.530 107.000 ;
        RECT 193.270 106.800 193.590 106.860 ;
        RECT 418.210 106.800 418.530 106.860 ;
      LAYER via ;
        RECT 193.300 106.800 193.560 107.060 ;
        RECT 418.240 106.800 418.500 107.060 ;
      LAYER met2 ;
        RECT 419.410 500.000 419.690 504.000 ;
        RECT 419.450 498.340 419.590 500.000 ;
        RECT 418.760 498.200 419.590 498.340 ;
        RECT 418.760 472.840 418.900 498.200 ;
        RECT 418.300 472.700 418.900 472.840 ;
        RECT 418.300 107.090 418.440 472.700 ;
        RECT 193.300 106.770 193.560 107.090 ;
        RECT 418.240 106.770 418.500 107.090 ;
        RECT 193.360 82.870 193.500 106.770 ;
        RECT 193.360 82.730 198.560 82.870 ;
        RECT 198.420 2.400 198.560 82.730 ;
        RECT 198.210 -4.800 198.770 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.920 499.700 459.240 499.760 ;
        RECT 457.170 499.560 459.240 499.700 ;
        RECT 457.170 496.640 457.310 499.560 ;
        RECT 458.920 499.500 459.240 499.560 ;
        RECT 467.890 496.640 468.210 496.700 ;
        RECT 457.170 496.500 468.210 496.640 ;
        RECT 467.890 496.440 468.210 496.500 ;
        RECT 467.890 488.480 468.210 488.540 ;
        RECT 669.370 488.480 669.690 488.540 ;
        RECT 467.890 488.340 669.690 488.480 ;
        RECT 467.890 488.280 468.210 488.340 ;
        RECT 669.370 488.280 669.690 488.340 ;
      LAYER via ;
        RECT 458.950 499.500 459.210 499.760 ;
        RECT 467.920 496.440 468.180 496.700 ;
        RECT 467.920 488.280 468.180 488.540 ;
        RECT 669.400 488.280 669.660 488.540 ;
      LAYER met2 ;
        RECT 458.970 500.000 459.250 504.000 ;
        RECT 459.010 499.790 459.150 500.000 ;
        RECT 458.950 499.470 459.210 499.790 ;
        RECT 467.920 496.410 468.180 496.730 ;
        RECT 467.980 488.570 468.120 496.410 ;
        RECT 467.920 488.250 468.180 488.570 ;
        RECT 669.400 488.250 669.660 488.570 ;
        RECT 669.460 82.870 669.600 488.250 ;
        RECT 669.460 82.730 673.280 82.870 ;
        RECT 673.140 2.400 673.280 82.730 ;
        RECT 672.930 -4.800 673.490 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 460.990 488.140 461.310 488.200 ;
        RECT 679.490 488.140 679.810 488.200 ;
        RECT 460.990 488.000 679.810 488.140 ;
        RECT 460.990 487.940 461.310 488.000 ;
        RECT 679.490 487.940 679.810 488.000 ;
        RECT 679.490 16.900 679.810 16.960 ;
        RECT 689.610 16.900 689.930 16.960 ;
        RECT 679.490 16.760 689.930 16.900 ;
        RECT 679.490 16.700 679.810 16.760 ;
        RECT 689.610 16.700 689.930 16.760 ;
      LAYER via ;
        RECT 461.020 487.940 461.280 488.200 ;
        RECT 679.520 487.940 679.780 488.200 ;
        RECT 679.520 16.700 679.780 16.960 ;
        RECT 689.640 16.700 689.900 16.960 ;
      LAYER met2 ;
        RECT 460.350 500.000 460.630 504.000 ;
        RECT 460.390 498.680 460.530 500.000 ;
        RECT 460.390 498.540 460.760 498.680 ;
        RECT 460.620 490.010 460.760 498.540 ;
        RECT 460.620 489.870 461.220 490.010 ;
        RECT 461.080 488.230 461.220 489.870 ;
        RECT 461.020 487.910 461.280 488.230 ;
        RECT 679.520 487.910 679.780 488.230 ;
        RECT 679.580 16.990 679.720 487.910 ;
        RECT 679.520 16.670 679.780 16.990 ;
        RECT 689.640 16.670 689.900 16.990 ;
        RECT 689.700 2.400 689.840 16.670 ;
        RECT 689.490 -4.800 690.050 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 389.230 500.380 389.550 500.440 ;
        RECT 389.230 500.240 421.430 500.380 ;
        RECT 389.230 500.180 389.550 500.240 ;
        RECT 421.290 499.760 421.430 500.240 ;
        RECT 421.200 499.500 421.520 499.760 ;
        RECT 272.390 487.120 272.710 487.180 ;
        RECT 389.230 487.120 389.550 487.180 ;
        RECT 272.390 486.980 389.550 487.120 ;
        RECT 272.390 486.920 272.710 486.980 ;
        RECT 389.230 486.920 389.550 486.980 ;
        RECT 220.410 19.620 220.730 19.680 ;
        RECT 272.390 19.620 272.710 19.680 ;
        RECT 220.410 19.480 272.710 19.620 ;
        RECT 220.410 19.420 220.730 19.480 ;
        RECT 272.390 19.420 272.710 19.480 ;
      LAYER via ;
        RECT 389.260 500.180 389.520 500.440 ;
        RECT 421.230 499.500 421.490 499.760 ;
        RECT 272.420 486.920 272.680 487.180 ;
        RECT 389.260 486.920 389.520 487.180 ;
        RECT 220.440 19.420 220.700 19.680 ;
        RECT 272.420 19.420 272.680 19.680 ;
      LAYER met2 ;
        RECT 389.260 500.150 389.520 500.470 ;
        RECT 389.320 487.210 389.460 500.150 ;
        RECT 421.250 500.000 421.530 504.000 ;
        RECT 421.290 499.790 421.430 500.000 ;
        RECT 421.230 499.470 421.490 499.790 ;
        RECT 272.420 486.890 272.680 487.210 ;
        RECT 389.260 486.890 389.520 487.210 ;
        RECT 272.480 19.710 272.620 486.890 ;
        RECT 220.440 19.390 220.700 19.710 ;
        RECT 272.420 19.390 272.680 19.710 ;
        RECT 220.500 2.400 220.640 19.390 ;
        RECT 220.290 -4.800 220.850 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.040 499.160 423.360 499.420 ;
        RECT 423.130 498.000 423.270 499.160 ;
        RECT 421.980 497.860 423.270 498.000 ;
        RECT 421.980 497.320 422.120 497.860 ;
        RECT 422.810 497.320 423.130 497.380 ;
        RECT 421.980 497.180 423.130 497.320 ;
        RECT 422.810 497.120 423.130 497.180 ;
        RECT 242.490 31.520 242.810 31.580 ;
        RECT 422.810 31.520 423.130 31.580 ;
        RECT 242.490 31.380 423.130 31.520 ;
        RECT 242.490 31.320 242.810 31.380 ;
        RECT 422.810 31.320 423.130 31.380 ;
      LAYER via ;
        RECT 423.070 499.160 423.330 499.420 ;
        RECT 422.840 497.120 423.100 497.380 ;
        RECT 242.520 31.320 242.780 31.580 ;
        RECT 422.840 31.320 423.100 31.580 ;
      LAYER met2 ;
        RECT 423.090 500.000 423.370 504.000 ;
        RECT 423.130 499.450 423.270 500.000 ;
        RECT 423.070 499.130 423.330 499.450 ;
        RECT 422.840 497.090 423.100 497.410 ;
        RECT 422.900 31.610 423.040 497.090 ;
        RECT 242.520 31.290 242.780 31.610 ;
        RECT 422.840 31.290 423.100 31.610 ;
        RECT 242.580 2.400 242.720 31.290 ;
        RECT 242.370 -4.800 242.930 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 313.790 488.140 314.110 488.200 ;
        RECT 421.430 488.140 421.750 488.200 ;
        RECT 313.790 488.000 421.750 488.140 ;
        RECT 313.790 487.940 314.110 488.000 ;
        RECT 421.430 487.940 421.750 488.000 ;
        RECT 259.050 19.960 259.370 20.020 ;
        RECT 313.790 19.960 314.110 20.020 ;
        RECT 259.050 19.820 314.110 19.960 ;
        RECT 259.050 19.760 259.370 19.820 ;
        RECT 313.790 19.760 314.110 19.820 ;
      LAYER via ;
        RECT 313.820 487.940 314.080 488.200 ;
        RECT 421.460 487.940 421.720 488.200 ;
        RECT 259.080 19.760 259.340 20.020 ;
        RECT 313.820 19.760 314.080 20.020 ;
      LAYER met2 ;
        RECT 424.470 500.000 424.750 504.000 ;
        RECT 424.510 498.965 424.650 500.000 ;
        RECT 421.450 498.595 421.730 498.965 ;
        RECT 424.440 498.595 424.720 498.965 ;
        RECT 421.520 488.230 421.660 498.595 ;
        RECT 313.820 487.910 314.080 488.230 ;
        RECT 421.460 487.910 421.720 488.230 ;
        RECT 313.880 20.050 314.020 487.910 ;
        RECT 259.080 19.730 259.340 20.050 ;
        RECT 313.820 19.730 314.080 20.050 ;
        RECT 259.140 2.400 259.280 19.730 ;
        RECT 258.930 -4.800 259.490 2.400 ;
      LAYER via2 ;
        RECT 421.450 498.640 421.730 498.920 ;
        RECT 424.440 498.640 424.720 498.920 ;
      LAYER met3 ;
        RECT 421.425 498.930 421.755 498.945 ;
        RECT 424.415 498.930 424.745 498.945 ;
        RECT 421.425 498.630 424.745 498.930 ;
        RECT 421.425 498.615 421.755 498.630 ;
        RECT 424.415 498.615 424.745 498.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 425.800 499.700 426.120 499.760 ;
        RECT 424.050 499.560 426.120 499.700 ;
        RECT 423.270 497.320 423.590 497.380 ;
        RECT 424.050 497.320 424.190 499.560 ;
        RECT 425.800 499.500 426.120 499.560 ;
        RECT 423.270 497.180 424.190 497.320 ;
        RECT 423.270 497.120 423.590 497.180 ;
        RECT 275.610 31.860 275.930 31.920 ;
        RECT 423.270 31.860 423.590 31.920 ;
        RECT 275.610 31.720 423.590 31.860 ;
        RECT 275.610 31.660 275.930 31.720 ;
        RECT 423.270 31.660 423.590 31.720 ;
      LAYER via ;
        RECT 423.300 497.120 423.560 497.380 ;
        RECT 425.830 499.500 426.090 499.760 ;
        RECT 275.640 31.660 275.900 31.920 ;
        RECT 423.300 31.660 423.560 31.920 ;
      LAYER met2 ;
        RECT 425.850 500.000 426.130 504.000 ;
        RECT 425.890 499.790 426.030 500.000 ;
        RECT 425.830 499.470 426.090 499.790 ;
        RECT 423.300 497.090 423.560 497.410 ;
        RECT 423.360 31.950 423.500 497.090 ;
        RECT 275.640 31.630 275.900 31.950 ;
        RECT 423.300 31.630 423.560 31.950 ;
        RECT 275.700 2.400 275.840 31.630 ;
        RECT 275.490 -4.800 276.050 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 355.190 485.080 355.510 485.140 ;
        RECT 427.410 485.080 427.730 485.140 ;
        RECT 355.190 484.940 427.730 485.080 ;
        RECT 355.190 484.880 355.510 484.940 ;
        RECT 427.410 484.880 427.730 484.940 ;
        RECT 292.170 19.620 292.490 19.680 ;
        RECT 355.190 19.620 355.510 19.680 ;
        RECT 292.170 19.480 355.510 19.620 ;
        RECT 292.170 19.420 292.490 19.480 ;
        RECT 355.190 19.420 355.510 19.480 ;
      LAYER via ;
        RECT 355.220 484.880 355.480 485.140 ;
        RECT 427.440 484.880 427.700 485.140 ;
        RECT 292.200 19.420 292.460 19.680 ;
        RECT 355.220 19.420 355.480 19.680 ;
      LAYER met2 ;
        RECT 427.230 500.000 427.510 504.000 ;
        RECT 427.270 498.850 427.410 500.000 ;
        RECT 427.270 498.710 427.640 498.850 ;
        RECT 427.500 485.170 427.640 498.710 ;
        RECT 355.220 484.850 355.480 485.170 ;
        RECT 427.440 484.850 427.700 485.170 ;
        RECT 355.280 19.710 355.420 484.850 ;
        RECT 292.200 19.390 292.460 19.710 ;
        RECT 355.220 19.390 355.480 19.710 ;
        RECT 292.260 2.400 292.400 19.390 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.250 472.840 429.570 472.900 ;
        RECT 431.550 472.840 431.870 472.900 ;
        RECT 429.250 472.700 431.870 472.840 ;
        RECT 429.250 472.640 429.570 472.700 ;
        RECT 431.550 472.640 431.870 472.700 ;
        RECT 308.730 38.320 309.050 38.380 ;
        RECT 431.550 38.320 431.870 38.380 ;
        RECT 308.730 38.180 431.870 38.320 ;
        RECT 308.730 38.120 309.050 38.180 ;
        RECT 431.550 38.120 431.870 38.180 ;
      LAYER via ;
        RECT 429.280 472.640 429.540 472.900 ;
        RECT 431.580 472.640 431.840 472.900 ;
        RECT 308.760 38.120 309.020 38.380 ;
        RECT 431.580 38.120 431.840 38.380 ;
      LAYER met2 ;
        RECT 428.610 500.000 428.890 504.000 ;
        RECT 428.650 499.645 428.790 500.000 ;
        RECT 428.580 499.275 428.860 499.645 ;
        RECT 428.810 498.595 429.090 498.965 ;
        RECT 428.880 498.170 429.020 498.595 ;
        RECT 428.880 498.030 429.480 498.170 ;
        RECT 429.340 472.930 429.480 498.030 ;
        RECT 429.280 472.610 429.540 472.930 ;
        RECT 431.580 472.610 431.840 472.930 ;
        RECT 431.640 38.410 431.780 472.610 ;
        RECT 308.760 38.090 309.020 38.410 ;
        RECT 431.580 38.090 431.840 38.410 ;
        RECT 308.820 2.400 308.960 38.090 ;
        RECT 308.610 -4.800 309.170 2.400 ;
      LAYER via2 ;
        RECT 428.580 499.320 428.860 499.600 ;
        RECT 428.810 498.640 429.090 498.920 ;
      LAYER met3 ;
        RECT 428.555 499.610 428.885 499.625 ;
        RECT 428.555 499.310 430.020 499.610 ;
        RECT 428.555 499.295 428.885 499.310 ;
        RECT 428.785 498.930 429.115 498.945 ;
        RECT 429.720 498.930 430.020 499.310 ;
        RECT 428.785 498.630 430.020 498.930 ;
        RECT 428.785 498.615 429.115 498.630 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 409.010 500.720 409.330 500.780 ;
        RECT 409.010 500.580 430.170 500.720 ;
        RECT 409.010 500.520 409.330 500.580 ;
        RECT 430.030 499.760 430.170 500.580 ;
        RECT 429.940 499.500 430.260 499.760 ;
        RECT 324.370 488.480 324.690 488.540 ;
        RECT 409.010 488.480 409.330 488.540 ;
        RECT 324.370 488.340 409.330 488.480 ;
        RECT 324.370 488.280 324.690 488.340 ;
        RECT 409.010 488.280 409.330 488.340 ;
      LAYER via ;
        RECT 409.040 500.520 409.300 500.780 ;
        RECT 429.970 499.500 430.230 499.760 ;
        RECT 324.400 488.280 324.660 488.540 ;
        RECT 409.040 488.280 409.300 488.540 ;
      LAYER met2 ;
        RECT 409.040 500.490 409.300 500.810 ;
        RECT 409.100 488.570 409.240 500.490 ;
        RECT 429.990 500.000 430.270 504.000 ;
        RECT 430.030 499.790 430.170 500.000 ;
        RECT 429.970 499.470 430.230 499.790 ;
        RECT 324.400 488.250 324.660 488.570 ;
        RECT 409.040 488.250 409.300 488.570 ;
        RECT 324.460 82.870 324.600 488.250 ;
        RECT 324.460 82.730 325.520 82.870 ;
        RECT 325.380 2.400 325.520 82.730 ;
        RECT 325.170 -4.800 325.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 416.140 498.820 416.460 499.080 ;
        RECT 416.230 498.680 416.370 498.820 ;
        RECT 416.230 498.540 417.060 498.680 ;
        RECT 416.920 497.720 417.060 498.540 ;
        RECT 416.830 497.460 417.150 497.720 ;
        RECT 416.830 490.860 417.150 490.920 ;
        RECT 419.590 490.860 419.910 490.920 ;
        RECT 416.830 490.720 419.910 490.860 ;
        RECT 416.830 490.660 417.150 490.720 ;
        RECT 419.590 490.660 419.910 490.720 ;
        RECT 158.770 424.560 159.090 424.620 ;
        RECT 419.590 424.560 419.910 424.620 ;
        RECT 158.770 424.420 419.910 424.560 ;
        RECT 158.770 424.360 159.090 424.420 ;
        RECT 419.590 424.360 419.910 424.420 ;
      LAYER via ;
        RECT 416.170 498.820 416.430 499.080 ;
        RECT 416.860 497.460 417.120 497.720 ;
        RECT 416.860 490.660 417.120 490.920 ;
        RECT 419.620 490.660 419.880 490.920 ;
        RECT 158.800 424.360 159.060 424.620 ;
        RECT 419.620 424.360 419.880 424.620 ;
      LAYER met2 ;
        RECT 416.190 500.000 416.470 504.000 ;
        RECT 416.230 499.110 416.370 500.000 ;
        RECT 416.170 498.790 416.430 499.110 ;
        RECT 416.860 497.430 417.120 497.750 ;
        RECT 416.920 490.950 417.060 497.430 ;
        RECT 416.860 490.630 417.120 490.950 ;
        RECT 419.620 490.630 419.880 490.950 ;
        RECT 419.680 424.650 419.820 490.630 ;
        RECT 158.800 424.330 159.060 424.650 ;
        RECT 419.620 424.330 419.880 424.650 ;
        RECT 158.860 82.870 159.000 424.330 ;
        RECT 158.860 82.730 159.920 82.870 ;
        RECT 159.780 2.400 159.920 82.730 ;
        RECT 159.570 -4.800 160.130 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.110 500.040 402.430 500.100 ;
        RECT 402.110 499.900 418.210 500.040 ;
        RECT 402.110 499.840 402.430 499.900 ;
        RECT 418.070 499.760 418.210 499.900 ;
        RECT 417.980 499.500 418.300 499.760 ;
        RECT 217.190 486.780 217.510 486.840 ;
        RECT 402.110 486.780 402.430 486.840 ;
        RECT 217.190 486.640 402.430 486.780 ;
        RECT 217.190 486.580 217.510 486.640 ;
        RECT 402.110 486.580 402.430 486.640 ;
        RECT 181.770 15.200 182.090 15.260 ;
        RECT 217.190 15.200 217.510 15.260 ;
        RECT 181.770 15.060 217.510 15.200 ;
        RECT 181.770 15.000 182.090 15.060 ;
        RECT 217.190 15.000 217.510 15.060 ;
      LAYER via ;
        RECT 402.140 499.840 402.400 500.100 ;
        RECT 418.010 499.500 418.270 499.760 ;
        RECT 217.220 486.580 217.480 486.840 ;
        RECT 402.140 486.580 402.400 486.840 ;
        RECT 181.800 15.000 182.060 15.260 ;
        RECT 217.220 15.000 217.480 15.260 ;
      LAYER met2 ;
        RECT 402.140 499.810 402.400 500.130 ;
        RECT 418.030 500.000 418.310 504.000 ;
        RECT 402.200 486.870 402.340 499.810 ;
        RECT 418.070 499.790 418.210 500.000 ;
        RECT 418.010 499.470 418.270 499.790 ;
        RECT 217.220 486.550 217.480 486.870 ;
        RECT 402.140 486.550 402.400 486.870 ;
        RECT 217.280 15.290 217.420 486.550 ;
        RECT 181.800 14.970 182.060 15.290 ;
        RECT 217.220 14.970 217.480 15.290 ;
        RECT 181.860 2.400 182.000 14.970 ;
        RECT 181.650 -4.800 182.210 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.170 438.160 200.490 438.220 ;
        RECT 420.050 438.160 420.370 438.220 ;
        RECT 200.170 438.020 420.370 438.160 ;
        RECT 200.170 437.960 200.490 438.020 ;
        RECT 420.050 437.960 420.370 438.020 ;
      LAYER via ;
        RECT 200.200 437.960 200.460 438.220 ;
        RECT 420.080 437.960 420.340 438.220 ;
      LAYER met2 ;
        RECT 419.870 500.000 420.150 504.000 ;
        RECT 419.910 498.850 420.050 500.000 ;
        RECT 419.910 498.710 420.280 498.850 ;
        RECT 420.140 438.250 420.280 498.710 ;
        RECT 200.200 437.930 200.460 438.250 ;
        RECT 420.080 437.930 420.340 438.250 ;
        RECT 200.260 82.870 200.400 437.930 ;
        RECT 200.260 82.730 204.080 82.870 ;
        RECT 203.940 2.400 204.080 82.730 ;
        RECT 203.730 -4.800 204.290 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.660 499.500 421.980 499.760 ;
        RECT 421.750 499.360 421.890 499.500 ;
        RECT 421.750 499.220 422.120 499.360 ;
        RECT 421.980 499.080 422.120 499.220 ;
        RECT 421.890 498.820 422.210 499.080 ;
        RECT 293.090 487.800 293.410 487.860 ;
        RECT 421.890 487.800 422.210 487.860 ;
        RECT 293.090 487.660 422.210 487.800 ;
        RECT 293.090 487.600 293.410 487.660 ;
        RECT 421.890 487.600 422.210 487.660 ;
        RECT 225.930 19.280 226.250 19.340 ;
        RECT 293.090 19.280 293.410 19.340 ;
        RECT 225.930 19.140 293.410 19.280 ;
        RECT 225.930 19.080 226.250 19.140 ;
        RECT 293.090 19.080 293.410 19.140 ;
      LAYER via ;
        RECT 421.690 499.500 421.950 499.760 ;
        RECT 421.920 498.820 422.180 499.080 ;
        RECT 293.120 487.600 293.380 487.860 ;
        RECT 421.920 487.600 422.180 487.860 ;
        RECT 225.960 19.080 226.220 19.340 ;
        RECT 293.120 19.080 293.380 19.340 ;
      LAYER met2 ;
        RECT 421.710 500.000 421.990 504.000 ;
        RECT 421.750 499.790 421.890 500.000 ;
        RECT 421.690 499.470 421.950 499.790 ;
        RECT 421.920 498.790 422.180 499.110 ;
        RECT 421.980 487.890 422.120 498.790 ;
        RECT 293.120 487.570 293.380 487.890 ;
        RECT 421.920 487.570 422.180 487.890 ;
        RECT 293.180 19.370 293.320 487.570 ;
        RECT 225.960 19.050 226.220 19.370 ;
        RECT 293.120 19.050 293.380 19.370 ;
        RECT 226.020 2.400 226.160 19.050 ;
        RECT 225.810 -4.800 226.370 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 413.840 499.160 414.160 499.420 ;
        RECT 413.930 498.340 414.070 499.160 ;
        RECT 414.530 498.340 414.850 498.400 ;
        RECT 413.930 498.200 414.850 498.340 ;
        RECT 414.530 498.140 414.850 498.200 ;
        RECT 414.530 472.160 414.850 472.220 ;
        RECT 417.290 472.160 417.610 472.220 ;
        RECT 414.530 472.020 417.610 472.160 ;
        RECT 414.530 471.960 414.850 472.020 ;
        RECT 417.290 471.960 417.610 472.020 ;
        RECT 132.090 37.980 132.410 38.040 ;
        RECT 417.290 37.980 417.610 38.040 ;
        RECT 132.090 37.840 417.610 37.980 ;
        RECT 132.090 37.780 132.410 37.840 ;
        RECT 417.290 37.780 417.610 37.840 ;
      LAYER via ;
        RECT 413.870 499.160 414.130 499.420 ;
        RECT 414.560 498.140 414.820 498.400 ;
        RECT 414.560 471.960 414.820 472.220 ;
        RECT 417.320 471.960 417.580 472.220 ;
        RECT 132.120 37.780 132.380 38.040 ;
        RECT 417.320 37.780 417.580 38.040 ;
      LAYER met2 ;
        RECT 413.890 500.000 414.170 504.000 ;
        RECT 413.930 499.450 414.070 500.000 ;
        RECT 413.870 499.130 414.130 499.450 ;
        RECT 414.560 498.110 414.820 498.430 ;
        RECT 414.620 472.250 414.760 498.110 ;
        RECT 414.560 471.930 414.820 472.250 ;
        RECT 417.320 471.930 417.580 472.250 ;
        RECT 417.380 38.070 417.520 471.930 ;
        RECT 132.120 37.750 132.380 38.070 ;
        RECT 417.320 37.750 417.580 38.070 ;
        RECT 132.180 2.400 132.320 37.750 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 155.090 486.440 155.410 486.500 ;
        RECT 414.070 486.440 414.390 486.500 ;
        RECT 155.090 486.300 414.390 486.440 ;
        RECT 155.090 486.240 155.410 486.300 ;
        RECT 414.070 486.240 414.390 486.300 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 155.090 17.580 155.410 17.640 ;
        RECT 137.610 17.440 155.410 17.580 ;
        RECT 137.610 17.380 137.930 17.440 ;
        RECT 155.090 17.380 155.410 17.440 ;
      LAYER via ;
        RECT 155.120 486.240 155.380 486.500 ;
        RECT 414.100 486.240 414.360 486.500 ;
        RECT 137.640 17.380 137.900 17.640 ;
        RECT 155.120 17.380 155.380 17.640 ;
      LAYER met2 ;
        RECT 414.350 500.000 414.630 504.000 ;
        RECT 414.390 498.850 414.530 500.000 ;
        RECT 414.160 498.710 414.530 498.850 ;
        RECT 414.160 486.530 414.300 498.710 ;
        RECT 155.120 486.210 155.380 486.530 ;
        RECT 414.100 486.210 414.360 486.530 ;
        RECT 155.180 17.670 155.320 486.210 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 155.120 17.350 155.380 17.670 ;
        RECT 137.700 2.400 137.840 17.350 ;
        RECT 137.490 -4.800 138.050 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 405.330 735.225 644.450 736.830 ;
        RECT 405.330 729.785 644.450 732.615 ;
        RECT 405.330 724.345 644.450 727.175 ;
        RECT 405.330 718.905 644.450 721.735 ;
        RECT 405.330 713.465 644.450 716.295 ;
        RECT 405.330 708.025 644.450 710.855 ;
        RECT 405.330 702.585 644.450 705.415 ;
        RECT 405.330 697.145 644.450 699.975 ;
        RECT 405.330 691.705 644.450 694.535 ;
        RECT 405.330 686.265 644.450 689.095 ;
        RECT 405.330 680.825 644.450 683.655 ;
        RECT 405.330 675.385 644.450 678.215 ;
        RECT 405.330 669.945 644.450 672.775 ;
        RECT 405.330 664.505 644.450 667.335 ;
        RECT 405.330 659.065 644.450 661.895 ;
        RECT 405.330 653.625 644.450 656.455 ;
        RECT 405.330 648.185 644.450 651.015 ;
        RECT 405.330 642.745 644.450 645.575 ;
        RECT 405.330 637.305 644.450 640.135 ;
        RECT 405.330 631.865 644.450 634.695 ;
        RECT 405.330 626.425 644.450 629.255 ;
        RECT 405.330 620.985 644.450 623.815 ;
        RECT 405.330 615.545 644.450 618.375 ;
        RECT 405.330 610.105 644.450 612.935 ;
        RECT 405.330 604.665 644.450 607.495 ;
        RECT 405.330 599.225 644.450 602.055 ;
        RECT 405.330 593.785 644.450 596.615 ;
        RECT 405.330 588.345 644.450 591.175 ;
        RECT 405.330 582.905 644.450 585.735 ;
        RECT 405.330 577.465 644.450 580.295 ;
        RECT 405.330 572.025 644.450 574.855 ;
        RECT 405.330 566.585 644.450 569.415 ;
        RECT 405.330 561.145 644.450 563.975 ;
        RECT 405.330 555.705 644.450 558.535 ;
        RECT 405.330 550.265 644.450 553.095 ;
        RECT 405.330 544.825 644.450 547.655 ;
        RECT 405.330 539.385 644.450 542.215 ;
        RECT 405.330 533.945 644.450 536.775 ;
        RECT 405.330 528.505 644.450 531.335 ;
        RECT 405.330 523.065 644.450 525.895 ;
        RECT 405.330 517.625 644.450 520.455 ;
        RECT 405.330 512.185 644.450 515.015 ;
      LAYER li1 ;
        RECT 405.520 510.795 644.260 736.725 ;
      LAYER met1 ;
        RECT 405.520 507.860 644.260 742.040 ;
      LAYER met2 ;
        RECT 412.980 745.720 424.190 746.570 ;
        RECT 425.030 745.720 425.570 746.570 ;
        RECT 426.410 745.720 426.950 746.570 ;
        RECT 427.790 745.720 428.330 746.570 ;
        RECT 429.170 745.720 429.710 746.570 ;
        RECT 430.550 745.720 431.090 746.570 ;
        RECT 431.930 745.720 432.470 746.570 ;
        RECT 433.310 745.720 433.850 746.570 ;
        RECT 434.690 745.720 435.230 746.570 ;
        RECT 436.070 745.720 436.610 746.570 ;
        RECT 437.450 745.720 437.990 746.570 ;
        RECT 438.830 745.720 439.370 746.570 ;
        RECT 440.210 745.720 440.750 746.570 ;
        RECT 441.590 745.720 442.130 746.570 ;
        RECT 442.970 745.720 443.510 746.570 ;
        RECT 444.350 745.720 444.890 746.570 ;
        RECT 445.730 745.720 446.270 746.570 ;
        RECT 447.110 745.720 447.650 746.570 ;
        RECT 448.490 745.720 449.030 746.570 ;
        RECT 449.870 745.720 450.410 746.570 ;
        RECT 451.250 745.720 451.790 746.570 ;
        RECT 452.630 745.720 453.170 746.570 ;
        RECT 454.010 745.720 454.550 746.570 ;
        RECT 455.390 745.720 455.930 746.570 ;
        RECT 456.770 745.720 457.310 746.570 ;
        RECT 458.150 745.720 458.690 746.570 ;
        RECT 459.530 745.720 460.070 746.570 ;
        RECT 460.910 745.720 461.450 746.570 ;
        RECT 462.290 745.720 462.830 746.570 ;
        RECT 463.670 745.720 464.210 746.570 ;
        RECT 465.050 745.720 465.590 746.570 ;
        RECT 466.430 745.720 466.970 746.570 ;
        RECT 467.810 745.720 468.350 746.570 ;
        RECT 469.190 745.720 469.730 746.570 ;
        RECT 470.570 745.720 471.110 746.570 ;
        RECT 471.950 745.720 472.490 746.570 ;
        RECT 473.330 745.720 473.870 746.570 ;
        RECT 474.710 745.720 475.250 746.570 ;
        RECT 476.090 745.720 476.630 746.570 ;
        RECT 477.470 745.720 478.010 746.570 ;
        RECT 478.850 745.720 479.390 746.570 ;
        RECT 480.230 745.720 480.770 746.570 ;
        RECT 481.610 745.720 482.150 746.570 ;
        RECT 482.990 745.720 483.530 746.570 ;
        RECT 484.370 745.720 484.910 746.570 ;
        RECT 485.750 745.720 486.290 746.570 ;
        RECT 487.130 745.720 487.670 746.570 ;
        RECT 488.510 745.720 489.050 746.570 ;
        RECT 489.890 745.720 490.430 746.570 ;
        RECT 491.270 745.720 491.810 746.570 ;
        RECT 492.650 745.720 493.190 746.570 ;
        RECT 494.030 745.720 494.570 746.570 ;
        RECT 495.410 745.720 495.950 746.570 ;
        RECT 496.790 745.720 497.330 746.570 ;
        RECT 498.170 745.720 498.710 746.570 ;
        RECT 499.550 745.720 500.090 746.570 ;
        RECT 500.930 745.720 501.470 746.570 ;
        RECT 502.310 745.720 502.850 746.570 ;
        RECT 503.690 745.720 504.230 746.570 ;
        RECT 505.070 745.720 505.610 746.570 ;
        RECT 506.450 745.720 506.990 746.570 ;
        RECT 507.830 745.720 508.370 746.570 ;
        RECT 509.210 745.720 509.750 746.570 ;
        RECT 510.590 745.720 511.130 746.570 ;
        RECT 511.970 745.720 512.510 746.570 ;
        RECT 513.350 745.720 513.890 746.570 ;
        RECT 514.730 745.720 515.270 746.570 ;
        RECT 516.110 745.720 516.650 746.570 ;
        RECT 517.490 745.720 518.030 746.570 ;
        RECT 518.870 745.720 519.410 746.570 ;
        RECT 520.250 745.720 520.790 746.570 ;
        RECT 521.630 745.720 522.170 746.570 ;
        RECT 523.010 745.720 523.550 746.570 ;
        RECT 524.390 745.720 524.930 746.570 ;
        RECT 525.770 745.720 526.310 746.570 ;
        RECT 527.150 745.720 527.690 746.570 ;
        RECT 528.530 745.720 529.070 746.570 ;
        RECT 529.910 745.720 530.450 746.570 ;
        RECT 531.290 745.720 531.830 746.570 ;
        RECT 532.670 745.720 533.210 746.570 ;
        RECT 534.050 745.720 534.590 746.570 ;
        RECT 535.430 745.720 535.970 746.570 ;
        RECT 536.810 745.720 537.350 746.570 ;
        RECT 538.190 745.720 538.730 746.570 ;
        RECT 539.570 745.720 540.110 746.570 ;
        RECT 540.950 745.720 541.490 746.570 ;
        RECT 542.330 745.720 542.870 746.570 ;
        RECT 543.710 745.720 544.250 746.570 ;
        RECT 545.090 745.720 545.630 746.570 ;
        RECT 546.470 745.720 547.010 746.570 ;
        RECT 547.850 745.720 548.390 746.570 ;
        RECT 549.230 745.720 549.770 746.570 ;
        RECT 550.610 745.720 551.150 746.570 ;
        RECT 551.990 745.720 552.530 746.570 ;
        RECT 553.370 745.720 553.910 746.570 ;
        RECT 554.750 745.720 555.290 746.570 ;
        RECT 556.130 745.720 556.670 746.570 ;
        RECT 557.510 745.720 558.050 746.570 ;
        RECT 558.890 745.720 559.430 746.570 ;
        RECT 560.270 745.720 560.810 746.570 ;
        RECT 561.650 745.720 562.190 746.570 ;
        RECT 563.030 745.720 563.570 746.570 ;
        RECT 564.410 745.720 564.950 746.570 ;
        RECT 565.790 745.720 566.330 746.570 ;
        RECT 567.170 745.720 567.710 746.570 ;
        RECT 568.550 745.720 569.090 746.570 ;
        RECT 569.930 745.720 570.470 746.570 ;
        RECT 571.310 745.720 571.850 746.570 ;
        RECT 572.690 745.720 573.230 746.570 ;
        RECT 574.070 745.720 574.610 746.570 ;
        RECT 575.450 745.720 575.990 746.570 ;
        RECT 576.830 745.720 577.370 746.570 ;
        RECT 578.210 745.720 578.750 746.570 ;
        RECT 579.590 745.720 580.130 746.570 ;
        RECT 580.970 745.720 581.510 746.570 ;
        RECT 582.350 745.720 582.890 746.570 ;
        RECT 583.730 745.720 584.270 746.570 ;
        RECT 585.110 745.720 585.650 746.570 ;
        RECT 586.490 745.720 587.030 746.570 ;
        RECT 587.870 745.720 588.410 746.570 ;
        RECT 589.250 745.720 589.790 746.570 ;
        RECT 590.630 745.720 591.170 746.570 ;
        RECT 592.010 745.720 592.550 746.570 ;
        RECT 593.390 745.720 593.930 746.570 ;
        RECT 594.770 745.720 595.310 746.570 ;
        RECT 596.150 745.720 596.690 746.570 ;
        RECT 597.530 745.720 598.070 746.570 ;
        RECT 598.910 745.720 599.450 746.570 ;
        RECT 600.290 745.720 600.830 746.570 ;
        RECT 601.670 745.720 602.210 746.570 ;
        RECT 603.050 745.720 603.590 746.570 ;
        RECT 604.430 745.720 604.970 746.570 ;
        RECT 605.810 745.720 606.350 746.570 ;
        RECT 607.190 745.720 607.730 746.570 ;
        RECT 608.570 745.720 609.110 746.570 ;
        RECT 609.950 745.720 610.490 746.570 ;
        RECT 611.330 745.720 611.870 746.570 ;
        RECT 612.710 745.720 613.250 746.570 ;
        RECT 614.090 745.720 614.630 746.570 ;
        RECT 615.470 745.720 616.010 746.570 ;
        RECT 616.850 745.720 617.390 746.570 ;
        RECT 618.230 745.720 618.770 746.570 ;
        RECT 619.610 745.720 620.150 746.570 ;
        RECT 620.990 745.720 621.530 746.570 ;
        RECT 622.370 745.720 622.910 746.570 ;
        RECT 623.750 745.720 624.290 746.570 ;
        RECT 625.130 745.720 636.800 746.570 ;
        RECT 412.980 504.280 636.800 745.720 ;
      LAYER met2 ;
        RECT 412.050 500.000 412.330 504.000 ;
      LAYER met3 ;
        RECT 421.050 510.715 614.755 741.905 ;
      LAYER met4 ;
        RECT 507.935 737.280 578.185 741.905 ;
        RECT 507.935 517.175 574.240 737.280 ;
        RECT 576.640 517.175 578.185 737.280 ;
  END
END user_project_wrapper
END LIBRARY

