magic
tech sky130B
magscale 1 2
timestamp 1664920552
<< metal1 >>
rect 74534 702992 74540 703044
rect 74592 703032 74598 703044
rect 75730 703032 75736 703044
rect 74592 703004 75736 703032
rect 74592 702992 74598 703004
rect 75730 702992 75736 703004
rect 75788 702992 75794 703044
rect 204254 702992 204260 703044
rect 204312 703032 204318 703044
rect 205450 703032 205456 703044
rect 204312 703004 205456 703032
rect 204312 702992 204318 703004
rect 205450 702992 205456 703004
rect 205508 702992 205514 703044
rect 333974 702992 333980 703044
rect 334032 703032 334038 703044
rect 335170 703032 335176 703044
rect 334032 703004 335176 703032
rect 334032 702992 334038 703004
rect 335170 702992 335176 703004
rect 335228 702992 335234 703044
rect 463694 702992 463700 703044
rect 463752 703032 463758 703044
rect 464890 703032 464896 703044
rect 463752 703004 464896 703032
rect 463752 702992 463758 703004
rect 464890 702992 464896 703004
rect 464948 702992 464954 703044
rect 97350 700748 97356 700800
rect 97408 700788 97414 700800
rect 109034 700788 109040 700800
rect 97408 700760 109040 700788
rect 97408 700748 97414 700760
rect 109034 700748 109040 700760
rect 109092 700748 109098 700800
rect 107654 700680 107660 700732
rect 107712 700720 107718 700732
rect 162210 700720 162216 700732
rect 107712 700692 162216 700720
rect 107712 700680 107718 700692
rect 162210 700680 162216 700692
rect 162268 700680 162274 700732
rect 32490 700612 32496 700664
rect 32548 700652 32554 700664
rect 110966 700652 110972 700664
rect 32548 700624 110972 700652
rect 32548 700612 32554 700624
rect 110966 700612 110972 700624
rect 111024 700612 111030 700664
rect 107746 700544 107752 700596
rect 107804 700584 107810 700596
rect 227070 700584 227076 700596
rect 107804 700556 227076 700584
rect 107804 700544 107810 700556
rect 227070 700544 227076 700556
rect 227128 700544 227134 700596
rect 106274 700476 106280 700528
rect 106332 700516 106338 700528
rect 291930 700516 291936 700528
rect 106332 700488 291936 700516
rect 106332 700476 106338 700488
rect 291930 700476 291936 700488
rect 291988 700476 291994 700528
rect 103514 700408 103520 700460
rect 103572 700448 103578 700460
rect 421650 700448 421656 700460
rect 103572 700420 421656 700448
rect 103572 700408 103578 700420
rect 421650 700408 421656 700420
rect 421708 700408 421714 700460
rect 102134 700340 102140 700392
rect 102192 700380 102198 700392
rect 486510 700380 486516 700392
rect 102192 700352 486516 700380
rect 102192 700340 102198 700352
rect 486510 700340 486516 700352
rect 486568 700340 486574 700392
rect 102226 700272 102232 700324
rect 102284 700312 102290 700324
rect 551370 700312 551376 700324
rect 102284 700284 551376 700312
rect 102284 700272 102290 700284
rect 551370 700272 551376 700284
rect 551428 700272 551434 700324
rect 100846 695512 100852 695564
rect 100904 695552 100910 695564
rect 580166 695552 580172 695564
rect 100904 695524 580172 695552
rect 100904 695512 100910 695524
rect 580166 695512 580172 695524
rect 580224 695512 580230 695564
rect 3418 694152 3424 694204
rect 3476 694192 3482 694204
rect 111242 694192 111248 694204
rect 3476 694164 111248 694192
rect 3476 694152 3482 694164
rect 111242 694152 111248 694164
rect 111300 694152 111306 694204
rect 101030 680348 101036 680400
rect 101088 680388 101094 680400
rect 580166 680388 580172 680400
rect 101088 680360 580172 680388
rect 101088 680348 101094 680360
rect 580166 680348 580172 680360
rect 580224 680348 580230 680400
rect 3418 677560 3424 677612
rect 3476 677600 3482 677612
rect 112162 677600 112168 677612
rect 3476 677572 112168 677600
rect 3476 677560 3482 677572
rect 112162 677560 112168 677572
rect 112220 677560 112226 677612
rect 100202 663756 100208 663808
rect 100260 663796 100266 663808
rect 580166 663796 580172 663808
rect 100260 663768 580172 663796
rect 100260 663756 100266 663768
rect 580166 663756 580172 663768
rect 580224 663756 580230 663808
rect 3418 661036 3424 661088
rect 3476 661076 3482 661088
rect 111886 661076 111892 661088
rect 3476 661048 111892 661076
rect 3476 661036 3482 661048
rect 111886 661036 111892 661048
rect 111944 661036 111950 661088
rect 99650 648592 99656 648644
rect 99708 648632 99714 648644
rect 580166 648632 580172 648644
rect 99708 648604 580172 648632
rect 99708 648592 99714 648604
rect 580166 648592 580172 648604
rect 580224 648592 580230 648644
rect 3234 644444 3240 644496
rect 3292 644484 3298 644496
rect 112346 644484 112352 644496
rect 3292 644456 112352 644484
rect 3292 644444 3298 644456
rect 112346 644444 112352 644456
rect 112404 644444 112410 644496
rect 99926 633428 99932 633480
rect 99984 633468 99990 633480
rect 580166 633468 580172 633480
rect 99984 633440 580172 633468
rect 99984 633428 99990 633440
rect 580166 633428 580172 633440
rect 580224 633428 580230 633480
rect 3418 627920 3424 627972
rect 3476 627960 3482 627972
rect 113358 627960 113364 627972
rect 3476 627932 113364 627960
rect 3476 627920 3482 627932
rect 113358 627920 113364 627932
rect 113416 627920 113422 627972
rect 99466 616836 99472 616888
rect 99524 616876 99530 616888
rect 580166 616876 580172 616888
rect 99524 616848 580172 616876
rect 99524 616836 99530 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 111058 610008 111064 610020
rect 3476 609980 111064 610008
rect 3476 609968 3482 609980
rect 111058 609968 111064 609980
rect 111116 609968 111122 610020
rect 98546 601672 98552 601724
rect 98604 601712 98610 601724
rect 580166 601712 580172 601724
rect 98604 601684 580172 601712
rect 98604 601672 98610 601684
rect 580166 601672 580172 601684
rect 580224 601672 580230 601724
rect 98270 586508 98276 586560
rect 98328 586548 98334 586560
rect 580902 586548 580908 586560
rect 98328 586520 580908 586548
rect 98328 586508 98334 586520
rect 580902 586508 580908 586520
rect 580960 586508 580966 586560
rect 3050 576852 3056 576904
rect 3108 576892 3114 576904
rect 114002 576892 114008 576904
rect 3108 576864 114008 576892
rect 3108 576852 3114 576864
rect 114002 576852 114008 576864
rect 114060 576852 114066 576904
rect 98362 569916 98368 569968
rect 98420 569956 98426 569968
rect 580166 569956 580172 569968
rect 98420 569928 580172 569956
rect 98420 569916 98426 569928
rect 580166 569916 580172 569928
rect 580224 569916 580230 569968
rect 3050 560260 3056 560312
rect 3108 560300 3114 560312
rect 112438 560300 112444 560312
rect 3108 560272 112444 560300
rect 3108 560260 3114 560272
rect 112438 560260 112444 560272
rect 112496 560260 112502 560312
rect 97442 554752 97448 554804
rect 97500 554792 97506 554804
rect 580166 554792 580172 554804
rect 97500 554764 580172 554792
rect 97500 554752 97506 554764
rect 580166 554752 580172 554764
rect 580224 554752 580230 554804
rect 96890 539588 96896 539640
rect 96948 539628 96954 539640
rect 580166 539628 580172 539640
rect 96948 539600 580172 539628
rect 96948 539588 96954 539600
rect 580166 539588 580172 539600
rect 580224 539588 580230 539640
rect 3602 527144 3608 527196
rect 3660 527184 3666 527196
rect 115106 527184 115112 527196
rect 3660 527156 115112 527184
rect 3660 527144 3666 527156
rect 115106 527144 115112 527156
rect 115164 527144 115170 527196
rect 97166 522996 97172 523048
rect 97224 523036 97230 523048
rect 580166 523036 580172 523048
rect 97224 523008 580172 523036
rect 97224 522996 97230 523008
rect 580166 522996 580172 523008
rect 580224 522996 580230 523048
rect 3326 510620 3332 510672
rect 3384 510660 3390 510672
rect 112530 510660 112536 510672
rect 3384 510632 112536 510660
rect 3384 510620 3390 510632
rect 112530 510620 112536 510632
rect 112588 510620 112594 510672
rect 95786 507832 95792 507884
rect 95844 507872 95850 507884
rect 580166 507872 580172 507884
rect 95844 507844 580172 507872
rect 95844 507832 95850 507844
rect 580166 507832 580172 507844
rect 580224 507832 580230 507884
rect 3326 494028 3332 494080
rect 3384 494068 3390 494080
rect 116486 494068 116492 494080
rect 3384 494040 116492 494068
rect 3384 494028 3390 494040
rect 116486 494028 116492 494040
rect 116544 494028 116550 494080
rect 96706 492668 96712 492720
rect 96764 492708 96770 492720
rect 580166 492708 580172 492720
rect 96764 492680 580172 492708
rect 96764 492668 96770 492680
rect 580166 492668 580172 492680
rect 580224 492668 580230 492720
rect 3142 476144 3148 476196
rect 3200 476184 3206 476196
rect 116762 476184 116768 476196
rect 3200 476156 116768 476184
rect 3200 476144 3206 476156
rect 116762 476144 116768 476156
rect 116820 476144 116826 476196
rect 95510 476076 95516 476128
rect 95568 476116 95574 476128
rect 580166 476116 580172 476128
rect 95568 476088 580172 476116
rect 95568 476076 95574 476088
rect 580166 476076 580172 476088
rect 580224 476076 580230 476128
rect 95326 460912 95332 460964
rect 95384 460952 95390 460964
rect 580166 460952 580172 460964
rect 95384 460924 580172 460952
rect 95384 460912 95390 460924
rect 580166 460912 580172 460924
rect 580224 460912 580230 460964
rect 3142 459552 3148 459604
rect 3200 459592 3206 459604
rect 113818 459592 113824 459604
rect 3200 459564 113824 459592
rect 3200 459552 3206 459564
rect 113818 459552 113824 459564
rect 113876 459552 113882 459604
rect 95602 445748 95608 445800
rect 95660 445788 95666 445800
rect 580166 445788 580172 445800
rect 95660 445760 580172 445788
rect 95660 445748 95666 445760
rect 580166 445748 580172 445760
rect 580224 445748 580230 445800
rect 3326 442960 3332 443012
rect 3384 443000 3390 443012
rect 117038 443000 117044 443012
rect 3384 442972 117044 443000
rect 3384 442960 3390 442972
rect 117038 442960 117044 442972
rect 117096 442960 117102 443012
rect 94682 429156 94688 429208
rect 94740 429196 94746 429208
rect 580166 429196 580172 429208
rect 94740 429168 580172 429196
rect 94740 429156 94746 429168
rect 580166 429156 580172 429168
rect 580224 429156 580230 429208
rect 3326 426436 3332 426488
rect 3384 426476 3390 426488
rect 117590 426476 117596 426488
rect 3384 426448 117596 426476
rect 3384 426436 3390 426448
rect 117590 426436 117596 426448
rect 117648 426436 117654 426488
rect 94130 413992 94136 414044
rect 94188 414032 94194 414044
rect 580166 414032 580172 414044
rect 94188 414004 580172 414032
rect 94188 413992 94194 414004
rect 580166 413992 580172 414004
rect 580224 413992 580230 414044
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 113910 409884 113916 409896
rect 3384 409856 113916 409884
rect 3384 409844 3390 409856
rect 113910 409844 113916 409856
rect 113968 409844 113974 409896
rect 94406 398828 94412 398880
rect 94464 398868 94470 398880
rect 580166 398868 580172 398880
rect 94464 398840 580172 398868
rect 94464 398828 94470 398840
rect 580166 398828 580172 398840
rect 580224 398828 580230 398880
rect 3602 393320 3608 393372
rect 3660 393360 3666 393372
rect 117866 393360 117872 393372
rect 3660 393332 117872 393360
rect 3660 393320 3666 393332
rect 117866 393320 117872 393332
rect 117924 393320 117930 393372
rect 93946 382236 93952 382288
rect 94004 382276 94010 382288
rect 580166 382276 580172 382288
rect 94004 382248 580172 382276
rect 94004 382236 94010 382248
rect 580166 382236 580172 382248
rect 580224 382236 580230 382288
rect 3326 376728 3332 376780
rect 3384 376768 3390 376780
rect 117958 376768 117964 376780
rect 3384 376740 117964 376768
rect 3384 376728 3390 376740
rect 117958 376728 117964 376740
rect 118016 376728 118022 376780
rect 92474 367072 92480 367124
rect 92532 367112 92538 367124
rect 580166 367112 580172 367124
rect 92532 367084 580172 367112
rect 92532 367072 92538 367084
rect 580166 367072 580172 367084
rect 580224 367072 580230 367124
rect 3326 360204 3332 360256
rect 3384 360244 3390 360256
rect 115198 360244 115204 360256
rect 3384 360216 115204 360244
rect 3384 360204 3390 360216
rect 115198 360204 115204 360216
rect 115256 360204 115262 360256
rect 92750 351908 92756 351960
rect 92808 351948 92814 351960
rect 580166 351948 580172 351960
rect 92808 351920 580172 351948
rect 92808 351908 92814 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 342252 3332 342304
rect 3384 342292 3390 342304
rect 119338 342292 119344 342304
rect 3384 342264 119344 342292
rect 3384 342252 3390 342264
rect 119338 342252 119344 342264
rect 119396 342252 119402 342304
rect 92842 335316 92848 335368
rect 92900 335356 92906 335368
rect 580166 335356 580172 335368
rect 92900 335328 580172 335356
rect 92900 335316 92906 335328
rect 580166 335316 580172 335328
rect 580224 335316 580230 335368
rect 3326 325660 3332 325712
rect 3384 325700 3390 325712
rect 118050 325700 118056 325712
rect 3384 325672 118056 325700
rect 3384 325660 3390 325672
rect 118050 325660 118056 325672
rect 118108 325660 118114 325712
rect 91094 320152 91100 320204
rect 91152 320192 91158 320204
rect 580166 320192 580172 320204
rect 91152 320164 580172 320192
rect 91152 320152 91158 320164
rect 580166 320152 580172 320164
rect 580224 320152 580230 320204
rect 3326 309136 3332 309188
rect 3384 309176 3390 309188
rect 119614 309176 119620 309188
rect 3384 309148 119620 309176
rect 3384 309136 3390 309148
rect 119614 309136 119620 309148
rect 119672 309136 119678 309188
rect 91370 304988 91376 305040
rect 91428 305028 91434 305040
rect 580166 305028 580172 305040
rect 91428 305000 580172 305028
rect 91428 304988 91434 305000
rect 580166 304988 580172 305000
rect 580224 304988 580230 305040
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 120626 292584 120632 292596
rect 3384 292556 120632 292584
rect 3384 292544 3390 292556
rect 120626 292544 120632 292556
rect 120684 292544 120690 292596
rect 91646 288396 91652 288448
rect 91704 288436 91710 288448
rect 580166 288436 580172 288448
rect 91704 288408 580172 288436
rect 91704 288396 91710 288408
rect 580166 288396 580172 288408
rect 580224 288396 580230 288448
rect 3326 276020 3332 276072
rect 3384 276060 3390 276072
rect 120718 276060 120724 276072
rect 3384 276032 120724 276060
rect 3384 276020 3390 276032
rect 120718 276020 120724 276032
rect 120776 276020 120782 276072
rect 89714 273232 89720 273284
rect 89772 273272 89778 273284
rect 580166 273272 580172 273284
rect 89772 273244 580172 273272
rect 89772 273232 89778 273244
rect 580166 273232 580172 273244
rect 580224 273232 580230 273284
rect 2958 259428 2964 259480
rect 3016 259468 3022 259480
rect 120442 259468 120448 259480
rect 3016 259440 120448 259468
rect 3016 259428 3022 259440
rect 120442 259428 120448 259440
rect 120500 259428 120506 259480
rect 91186 258068 91192 258120
rect 91244 258108 91250 258120
rect 580902 258108 580908 258120
rect 91244 258080 580908 258108
rect 91244 258068 91250 258080
rect 580902 258068 580908 258080
rect 580960 258068 580966 258120
rect 3326 242904 3332 242956
rect 3384 242944 3390 242956
rect 120350 242944 120356 242956
rect 3384 242916 120356 242944
rect 3384 242904 3390 242916
rect 120350 242904 120356 242916
rect 120408 242904 120414 242956
rect 89990 241476 89996 241528
rect 90048 241516 90054 241528
rect 580166 241516 580172 241528
rect 90048 241488 580172 241516
rect 90048 241476 90054 241488
rect 580166 241476 580172 241488
rect 580224 241476 580230 241528
rect 3326 226380 3332 226432
rect 3384 226420 3390 226432
rect 118142 226420 118148 226432
rect 3384 226392 118148 226420
rect 3384 226380 3390 226392
rect 118142 226380 118148 226392
rect 118200 226380 118206 226432
rect 89806 226312 89812 226364
rect 89864 226352 89870 226364
rect 580166 226352 580172 226364
rect 89864 226324 580172 226352
rect 89864 226312 89870 226324
rect 580166 226312 580172 226324
rect 580224 226312 580230 226364
rect 90082 211148 90088 211200
rect 90140 211188 90146 211200
rect 580166 211188 580172 211200
rect 90140 211160 580172 211188
rect 90140 211148 90146 211160
rect 580166 211148 580172 211160
rect 580224 211148 580230 211200
rect 3326 209788 3332 209840
rect 3384 209828 3390 209840
rect 116578 209828 116584 209840
rect 3384 209800 116584 209828
rect 3384 209788 3390 209800
rect 116578 209788 116584 209800
rect 116636 209788 116642 209840
rect 88334 194556 88340 194608
rect 88392 194596 88398 194608
rect 580166 194596 580172 194608
rect 88392 194568 580172 194596
rect 88392 194556 88398 194568
rect 580166 194556 580172 194568
rect 580224 194556 580230 194608
rect 3326 191836 3332 191888
rect 3384 191876 3390 191888
rect 121730 191876 121736 191888
rect 3384 191848 121736 191876
rect 3384 191836 3390 191848
rect 121730 191836 121736 191848
rect 121788 191836 121794 191888
rect 88610 179392 88616 179444
rect 88668 179432 88674 179444
rect 580166 179432 580172 179444
rect 88668 179404 580172 179432
rect 88668 179392 88674 179404
rect 580166 179392 580172 179404
rect 580224 179392 580230 179444
rect 3050 175244 3056 175296
rect 3108 175284 3114 175296
rect 122006 175284 122012 175296
rect 3108 175256 122012 175284
rect 3108 175244 3114 175256
rect 122006 175244 122012 175256
rect 122064 175244 122070 175296
rect 88886 164228 88892 164280
rect 88944 164268 88950 164280
rect 580166 164268 580172 164280
rect 88944 164240 580172 164268
rect 88944 164228 88950 164240
rect 580166 164228 580172 164240
rect 580224 164228 580230 164280
rect 88334 160216 88340 160268
rect 88392 160256 88398 160268
rect 89438 160256 89444 160268
rect 88392 160228 89444 160256
rect 88392 160216 88398 160228
rect 89438 160216 89444 160228
rect 89496 160216 89502 160268
rect 92750 159196 92756 159248
rect 92808 159236 92814 159248
rect 93302 159236 93308 159248
rect 92808 159208 93308 159236
rect 92808 159196 92814 159208
rect 93302 159196 93308 159208
rect 93360 159196 93366 159248
rect 107654 158856 107660 158908
rect 107712 158896 107718 158908
rect 108758 158896 108764 158908
rect 107712 158868 108764 158896
rect 107712 158856 107718 158868
rect 108758 158856 108764 158868
rect 108816 158856 108822 158908
rect 3142 158720 3148 158772
rect 3200 158760 3206 158772
rect 116486 158760 116492 158772
rect 3200 158732 116492 158760
rect 3200 158720 3206 158732
rect 116486 158720 116492 158732
rect 116544 158720 116550 158772
rect 102134 158244 102140 158296
rect 102192 158284 102198 158296
rect 103238 158284 103244 158296
rect 102192 158256 103244 158284
rect 102192 158244 102198 158256
rect 103238 158244 103244 158256
rect 103296 158244 103302 158296
rect 108482 157020 108488 157072
rect 108540 157060 108546 157072
rect 139394 157060 139400 157072
rect 108540 157032 139400 157060
rect 108540 157020 108546 157032
rect 139394 157020 139400 157032
rect 139452 157020 139458 157072
rect 74534 156952 74540 157004
rect 74592 156992 74598 157004
rect 109678 156992 109684 157004
rect 74592 156964 109684 156992
rect 74592 156952 74598 156964
rect 109678 156952 109684 156964
rect 109736 156952 109742 157004
rect 107378 156884 107384 156936
rect 107436 156924 107442 156936
rect 204254 156924 204260 156936
rect 107436 156896 204260 156924
rect 107436 156884 107442 156896
rect 204254 156884 204260 156896
rect 204312 156884 204318 156936
rect 9674 156816 9680 156868
rect 9732 156856 9738 156868
rect 110690 156856 110696 156868
rect 9732 156828 110696 156856
rect 9732 156816 9738 156828
rect 110690 156816 110696 156828
rect 110748 156816 110754 156868
rect 120350 156816 120356 156868
rect 120408 156856 120414 156868
rect 120902 156856 120908 156868
rect 120408 156828 120908 156856
rect 120408 156816 120414 156828
rect 120902 156816 120908 156828
rect 120960 156816 120966 156868
rect 106366 156748 106372 156800
rect 106424 156788 106430 156800
rect 269114 156788 269120 156800
rect 106424 156760 269120 156788
rect 106424 156748 106430 156760
rect 269114 156748 269120 156760
rect 269172 156748 269178 156800
rect 105078 156680 105084 156732
rect 105136 156720 105142 156732
rect 333974 156720 333980 156732
rect 105136 156692 333980 156720
rect 105136 156680 105142 156692
rect 333974 156680 333980 156692
rect 334032 156680 334038 156732
rect 105446 156612 105452 156664
rect 105504 156652 105510 156664
rect 356054 156652 356060 156664
rect 105504 156624 356060 156652
rect 105504 156612 105510 156624
rect 356054 156612 356060 156624
rect 356112 156612 356118 156664
rect 120350 156544 120356 156596
rect 120408 156584 120414 156596
rect 120626 156584 120632 156596
rect 120408 156556 120632 156584
rect 120408 156544 120414 156556
rect 120626 156544 120632 156556
rect 120684 156544 120690 156596
rect 113910 155864 113916 155916
rect 113968 155904 113974 155916
rect 117498 155904 117504 155916
rect 113968 155876 117504 155904
rect 113968 155864 113974 155876
rect 117498 155864 117504 155876
rect 117556 155864 117562 155916
rect 118050 155864 118056 155916
rect 118108 155904 118114 155916
rect 119798 155904 119804 155916
rect 118108 155876 119804 155904
rect 118108 155864 118114 155876
rect 119798 155864 119804 155876
rect 119856 155864 119862 155916
rect 108206 155592 108212 155644
rect 108264 155632 108270 155644
rect 183554 155632 183560 155644
rect 108264 155604 183560 155632
rect 108264 155592 108270 155604
rect 183554 155592 183560 155604
rect 183612 155592 183618 155644
rect 3418 155524 3424 155576
rect 3476 155564 3482 155576
rect 113726 155564 113732 155576
rect 3476 155536 113732 155564
rect 3476 155524 3482 155536
rect 113726 155524 113732 155536
rect 113784 155524 113790 155576
rect 3510 155456 3516 155508
rect 3568 155496 3574 155508
rect 114922 155496 114928 155508
rect 3568 155468 114928 155496
rect 3568 155456 3574 155468
rect 114922 155456 114928 155468
rect 114980 155456 114986 155508
rect 107102 155388 107108 155440
rect 107160 155428 107166 155440
rect 248414 155428 248420 155440
rect 107160 155400 248420 155428
rect 107160 155388 107166 155400
rect 248414 155388 248420 155400
rect 248472 155388 248478 155440
rect 104066 155320 104072 155372
rect 104124 155360 104130 155372
rect 398834 155360 398840 155372
rect 104124 155332 398840 155360
rect 104124 155320 104130 155332
rect 398834 155320 398840 155332
rect 398892 155320 398898 155372
rect 102962 155252 102968 155304
rect 103020 155292 103026 155304
rect 463694 155292 463700 155304
rect 103020 155264 463700 155292
rect 103020 155252 103026 155264
rect 463694 155252 463700 155264
rect 463752 155252 463758 155304
rect 101858 155184 101864 155236
rect 101916 155224 101922 155236
rect 528554 155224 528560 155236
rect 101916 155196 528560 155224
rect 101916 155184 101922 155196
rect 528554 155184 528560 155196
rect 528612 155184 528618 155236
rect 117958 154504 117964 154556
rect 118016 154544 118022 154556
rect 118694 154544 118700 154556
rect 118016 154516 118700 154544
rect 118016 154504 118022 154516
rect 118694 154504 118700 154516
rect 118752 154504 118758 154556
rect 109586 154232 109592 154284
rect 109644 154272 109650 154284
rect 118786 154272 118792 154284
rect 109644 154244 118792 154272
rect 109644 154232 109650 154244
rect 118786 154232 118792 154244
rect 118844 154232 118850 154284
rect 53834 154164 53840 154216
rect 53892 154204 53898 154216
rect 110414 154204 110420 154216
rect 53892 154176 110420 154204
rect 53892 154164 53898 154176
rect 110414 154164 110420 154176
rect 110472 154164 110478 154216
rect 106182 154096 106188 154148
rect 106240 154136 106246 154148
rect 313274 154136 313280 154148
rect 106240 154108 313280 154136
rect 106240 154096 106246 154108
rect 313274 154096 313280 154108
rect 313332 154096 313338 154148
rect 104986 154028 104992 154080
rect 105044 154068 105050 154080
rect 378134 154068 378140 154080
rect 105044 154040 378140 154068
rect 105044 154028 105050 154040
rect 378134 154028 378140 154040
rect 378192 154028 378198 154080
rect 103974 153960 103980 154012
rect 104032 154000 104038 154012
rect 442994 154000 443000 154012
rect 104032 153972 443000 154000
rect 104032 153960 104038 153972
rect 442994 153960 443000 153972
rect 443052 153960 443058 154012
rect 102870 153892 102876 153944
rect 102928 153932 102934 153944
rect 507854 153932 507860 153944
rect 102928 153904 507860 153932
rect 102928 153892 102934 153904
rect 507854 153892 507860 153904
rect 507912 153892 507918 153944
rect 101766 153824 101772 153876
rect 101824 153864 101830 153876
rect 572714 153864 572720 153876
rect 101824 153836 572720 153864
rect 101824 153824 101830 153836
rect 572714 153824 572720 153836
rect 572772 153824 572778 153876
rect 89990 153280 89996 153332
rect 90048 153320 90054 153332
rect 90542 153320 90548 153332
rect 90048 153292 90548 153320
rect 90048 153280 90054 153292
rect 90542 153280 90548 153292
rect 90600 153280 90606 153332
rect 91370 153280 91376 153332
rect 91428 153320 91434 153332
rect 92198 153320 92204 153332
rect 91428 153292 92204 153320
rect 91428 153280 91434 153292
rect 92198 153280 92204 153292
rect 92256 153280 92262 153332
rect 92474 153280 92480 153332
rect 92532 153320 92538 153332
rect 93026 153320 93032 153332
rect 92532 153292 93032 153320
rect 92532 153280 92538 153292
rect 93026 153280 93032 153292
rect 93084 153280 93090 153332
rect 95510 153280 95516 153332
rect 95568 153320 95574 153332
rect 96062 153320 96068 153332
rect 95568 153292 96068 153320
rect 95568 153280 95574 153292
rect 96062 153280 96068 153292
rect 96120 153280 96126 153332
rect 96890 153280 96896 153332
rect 96948 153320 96954 153332
rect 97718 153320 97724 153332
rect 96948 153292 97724 153320
rect 96948 153280 96954 153292
rect 97718 153280 97724 153292
rect 97776 153280 97782 153332
rect 98270 153280 98276 153332
rect 98328 153320 98334 153332
rect 98822 153320 98828 153332
rect 98328 153292 98828 153320
rect 98328 153280 98334 153292
rect 98822 153280 98828 153292
rect 98880 153280 98886 153332
rect 89714 153212 89720 153264
rect 89772 153252 89778 153264
rect 90818 153252 90824 153264
rect 89772 153224 90824 153252
rect 89772 153212 89778 153224
rect 90818 153212 90824 153224
rect 90876 153212 90882 153264
rect 91094 153212 91100 153264
rect 91152 153252 91158 153264
rect 91922 153252 91928 153264
rect 91152 153224 91928 153252
rect 91152 153212 91158 153224
rect 91922 153212 91928 153224
rect 91980 153212 91986 153264
rect 111058 153144 111064 153196
rect 111116 153184 111122 153196
rect 112898 153184 112904 153196
rect 111116 153156 112904 153184
rect 111116 153144 111122 153156
rect 112898 153144 112904 153156
rect 112956 153144 112962 153196
rect 113818 153144 113824 153196
rect 113876 153184 113882 153196
rect 116302 153184 116308 153196
rect 113876 153156 116308 153184
rect 113876 153144 113882 153156
rect 116302 153144 116308 153156
rect 116360 153144 116366 153196
rect 118142 153144 118148 153196
rect 118200 153184 118206 153196
rect 121454 153184 121460 153196
rect 118200 153156 121460 153184
rect 118200 153144 118206 153156
rect 121454 153144 121460 153156
rect 121512 153144 121518 153196
rect 115198 153076 115204 153128
rect 115256 153116 115262 153128
rect 118418 153116 118424 153128
rect 115256 153088 118424 153116
rect 115256 153076 115262 153088
rect 118418 153076 118424 153088
rect 118476 153076 118482 153128
rect 116578 153008 116584 153060
rect 116636 153048 116642 153060
rect 121178 153048 121184 153060
rect 116636 153020 121184 153048
rect 116636 153008 116642 153020
rect 121178 153008 121184 153020
rect 121236 153008 121242 153060
rect 116486 152940 116492 152992
rect 116544 152980 116550 152992
rect 122006 152980 122012 152992
rect 116544 152952 122012 152980
rect 116544 152940 116550 152952
rect 122006 152940 122012 152952
rect 122064 152940 122070 152992
rect 109310 152872 109316 152924
rect 109368 152912 109374 152924
rect 128722 152912 128728 152924
rect 109368 152884 128728 152912
rect 109368 152872 109374 152884
rect 128722 152872 128728 152884
rect 128780 152872 128786 152924
rect 123110 152844 123116 152856
rect 117884 152816 123116 152844
rect 7558 152668 7564 152720
rect 7616 152708 7622 152720
rect 117884 152708 117912 152816
rect 123110 152804 123116 152816
rect 123168 152804 123174 152856
rect 122834 152708 122840 152720
rect 7616 152680 117912 152708
rect 118160 152680 122840 152708
rect 7616 152668 7622 152680
rect 81894 152532 81900 152584
rect 81952 152572 81958 152584
rect 95786 152572 95792 152584
rect 81952 152544 95792 152572
rect 81952 152532 81958 152544
rect 95786 152532 95792 152544
rect 95844 152532 95850 152584
rect 80882 152464 80888 152516
rect 80940 152504 80946 152516
rect 94682 152504 94688 152516
rect 80940 152476 94688 152504
rect 80940 152464 80946 152476
rect 94682 152464 94688 152476
rect 94740 152464 94746 152516
rect 114830 152464 114836 152516
rect 114888 152504 114894 152516
rect 118050 152504 118056 152516
rect 114888 152476 118056 152504
rect 114888 152464 114894 152476
rect 118050 152464 118056 152476
rect 118108 152464 118114 152516
rect 4798 152396 4804 152448
rect 4856 152436 4862 152448
rect 118160 152436 118188 152680
rect 122834 152668 122840 152680
rect 122892 152668 122898 152720
rect 4856 152408 118188 152436
rect 4856 152396 4862 152408
rect 3786 152328 3792 152380
rect 3844 152368 3850 152380
rect 123938 152368 123944 152380
rect 3844 152340 123944 152368
rect 3844 152328 3850 152340
rect 123938 152328 123944 152340
rect 123996 152328 124002 152380
rect 82354 152260 82360 152312
rect 82412 152300 82418 152312
rect 101306 152300 101312 152312
rect 82412 152272 101312 152300
rect 82412 152260 82418 152272
rect 101306 152260 101312 152272
rect 101364 152260 101370 152312
rect 115842 152260 115848 152312
rect 115900 152300 115906 152312
rect 127986 152300 127992 152312
rect 115900 152272 127992 152300
rect 115900 152260 115906 152272
rect 127986 152260 127992 152272
rect 128044 152260 128050 152312
rect 82170 152192 82176 152244
rect 82228 152232 82234 152244
rect 96890 152232 96896 152244
rect 82228 152204 96896 152232
rect 82228 152192 82234 152204
rect 96890 152192 96896 152204
rect 96948 152192 96954 152244
rect 108114 152192 108120 152244
rect 108172 152232 108178 152244
rect 108172 152204 118004 152232
rect 108172 152192 108178 152204
rect 81710 152124 81716 152176
rect 81768 152164 81774 152176
rect 99098 152164 99104 152176
rect 81768 152136 99104 152164
rect 81768 152124 81774 152136
rect 99098 152124 99104 152136
rect 99156 152124 99162 152176
rect 111426 152124 111432 152176
rect 111484 152164 111490 152176
rect 117774 152164 117780 152176
rect 111484 152136 117780 152164
rect 111484 152124 111490 152136
rect 117774 152124 117780 152136
rect 117832 152124 117838 152176
rect 117976 152164 118004 152204
rect 118050 152192 118056 152244
rect 118108 152232 118114 152244
rect 128538 152232 128544 152244
rect 118108 152204 128544 152232
rect 118108 152192 118114 152204
rect 128538 152192 128544 152204
rect 128596 152192 128602 152244
rect 128446 152164 128452 152176
rect 117976 152136 128452 152164
rect 128446 152124 128452 152136
rect 128504 152124 128510 152176
rect 81434 152056 81440 152108
rect 81492 152096 81498 152108
rect 100202 152096 100208 152108
rect 81492 152068 100208 152096
rect 81492 152056 81498 152068
rect 100202 152056 100208 152068
rect 100260 152056 100266 152108
rect 104802 152056 104808 152108
rect 104860 152096 104866 152108
rect 128354 152096 128360 152108
rect 104860 152068 128360 152096
rect 104860 152056 104866 152068
rect 128354 152056 128360 152068
rect 128412 152056 128418 152108
rect 85850 151988 85856 152040
rect 85908 152028 85914 152040
rect 95234 152028 95240 152040
rect 85908 152000 95240 152028
rect 85908 151988 85914 152000
rect 95234 151988 95240 152000
rect 95292 151988 95298 152040
rect 103790 151988 103796 152040
rect 103848 152028 103854 152040
rect 128814 152028 128820 152040
rect 103848 152000 128820 152028
rect 103848 151988 103854 152000
rect 128814 151988 128820 152000
rect 128872 151988 128878 152040
rect 113634 151920 113640 151972
rect 113692 151960 113698 151972
rect 128906 151960 128912 151972
rect 113692 151932 128912 151960
rect 113692 151920 113698 151932
rect 128906 151920 128912 151932
rect 128964 151920 128970 151972
rect 112438 151852 112444 151904
rect 112496 151892 112502 151904
rect 114002 151892 114008 151904
rect 112496 151864 114008 151892
rect 112496 151852 112502 151864
rect 114002 151852 114008 151864
rect 114060 151852 114066 151904
rect 117774 151852 117780 151904
rect 117832 151892 117838 151904
rect 128630 151892 128636 151904
rect 117832 151864 128636 151892
rect 117832 151852 117838 151864
rect 128630 151852 128636 151864
rect 128688 151852 128694 151904
rect 82262 151784 82268 151836
rect 82320 151824 82326 151836
rect 98178 151824 98184 151836
rect 82320 151796 98184 151824
rect 82320 151784 82326 151796
rect 98178 151784 98184 151796
rect 98236 151784 98242 151836
rect 112530 151784 112536 151836
rect 112588 151824 112594 151836
rect 115014 151824 115020 151836
rect 112588 151796 115020 151824
rect 112588 151784 112594 151796
rect 115014 151784 115020 151796
rect 115072 151784 115078 151836
rect 116946 151784 116952 151836
rect 117004 151824 117010 151836
rect 128170 151824 128176 151836
rect 117004 151796 119200 151824
rect 117004 151784 117010 151796
rect 119172 151756 119200 151796
rect 120736 151796 128176 151824
rect 120736 151756 120764 151796
rect 128170 151784 128176 151796
rect 128228 151784 128234 151836
rect 119172 151728 120764 151756
rect 3510 151104 3516 151156
rect 3568 151144 3574 151156
rect 97994 151144 98000 151156
rect 3568 151116 98000 151144
rect 3568 151104 3574 151116
rect 97994 151104 98000 151116
rect 98052 151104 98058 151156
rect 95234 151036 95240 151088
rect 95292 151076 95298 151088
rect 580350 151076 580356 151088
rect 95292 151048 580356 151076
rect 95292 151036 95298 151048
rect 580350 151036 580356 151048
rect 580408 151036 580414 151088
rect 87782 150764 87788 150816
rect 87840 150804 87846 150816
rect 128998 150804 129004 150816
rect 87840 150776 129004 150804
rect 87840 150764 87846 150776
rect 128998 150764 129004 150776
rect 129056 150764 129062 150816
rect 3878 150696 3884 150748
rect 3936 150736 3942 150748
rect 123386 150736 123392 150748
rect 3936 150708 123392 150736
rect 3936 150696 3942 150708
rect 123386 150696 123392 150708
rect 123444 150696 123450 150748
rect 3694 150628 3700 150680
rect 3752 150668 3758 150680
rect 123662 150668 123668 150680
rect 3752 150640 123668 150668
rect 3752 150628 3758 150640
rect 123662 150628 123668 150640
rect 123720 150628 123726 150680
rect 3602 150560 3608 150612
rect 3660 150600 3666 150612
rect 124214 150600 124220 150612
rect 3660 150572 124220 150600
rect 3660 150560 3666 150572
rect 124214 150560 124220 150572
rect 124272 150560 124278 150612
rect 3234 150492 3240 150544
rect 3292 150532 3298 150544
rect 124490 150532 124496 150544
rect 3292 150504 124496 150532
rect 3292 150492 3298 150504
rect 124490 150492 124496 150504
rect 124548 150492 124554 150544
rect 88518 150424 88524 150476
rect 88576 150464 88582 150476
rect 580166 150464 580172 150476
rect 88576 150436 580172 150464
rect 88576 150424 88582 150436
rect 580166 150424 580172 150436
rect 580224 150424 580230 150476
rect 80974 150152 80980 150204
rect 81032 150192 81038 150204
rect 91508 150192 91514 150204
rect 81032 150164 91514 150192
rect 81032 150152 81038 150164
rect 91508 150152 91514 150164
rect 91566 150152 91572 150204
rect 81342 149948 81348 150000
rect 81400 149988 81406 150000
rect 81400 149960 89484 149988
rect 81400 149948 81406 149960
rect 81158 149880 81164 149932
rect 81216 149920 81222 149932
rect 81216 149892 89392 149920
rect 81216 149880 81222 149892
rect 81066 149744 81072 149796
rect 81124 149784 81130 149796
rect 89364 149784 89392 149892
rect 89456 149852 89484 149960
rect 93578 149852 93584 149864
rect 89456 149824 93584 149852
rect 93578 149812 93584 149824
rect 93636 149812 93642 149864
rect 112346 149812 112352 149864
rect 112404 149852 112410 149864
rect 112622 149852 112628 149864
rect 112404 149824 112628 149852
rect 112404 149812 112410 149824
rect 112622 149812 112628 149824
rect 112680 149812 112686 149864
rect 90266 149784 90272 149796
rect 81124 149756 89300 149784
rect 89364 149756 90272 149784
rect 81124 149744 81130 149756
rect 81250 149676 81256 149728
rect 81308 149716 81314 149728
rect 89162 149716 89168 149728
rect 81308 149688 89168 149716
rect 81308 149676 81314 149688
rect 89162 149676 89168 149688
rect 89220 149676 89226 149728
rect 89272 149716 89300 149756
rect 90266 149744 90272 149756
rect 90324 149744 90330 149796
rect 92474 149716 92480 149728
rect 89272 149688 92480 149716
rect 92474 149676 92480 149688
rect 92532 149676 92538 149728
rect 85298 149608 85304 149660
rect 85356 149648 85362 149660
rect 89438 149648 89444 149660
rect 85356 149620 89444 149648
rect 85356 149608 85362 149620
rect 89438 149608 89444 149620
rect 89496 149608 89502 149660
rect 91646 149608 91652 149660
rect 91704 149648 91710 149660
rect 91704 149620 99374 149648
rect 91704 149608 91710 149620
rect 81802 149540 81808 149592
rect 81860 149580 81866 149592
rect 86954 149580 86960 149592
rect 81860 149552 86960 149580
rect 81860 149540 81866 149552
rect 86954 149540 86960 149552
rect 87012 149540 87018 149592
rect 91922 149540 91928 149592
rect 91980 149580 91986 149592
rect 91980 149552 96614 149580
rect 91980 149540 91986 149552
rect 81986 149472 81992 149524
rect 82044 149512 82050 149524
rect 85850 149512 85856 149524
rect 82044 149484 85856 149512
rect 82044 149472 82050 149484
rect 85850 149472 85856 149484
rect 85908 149472 85914 149524
rect 85960 149484 86540 149512
rect 82078 149404 82084 149456
rect 82136 149444 82142 149456
rect 84562 149444 84568 149456
rect 82136 149416 84568 149444
rect 82136 149404 82142 149416
rect 84562 149404 84568 149416
rect 84620 149404 84626 149456
rect 3418 149336 3424 149388
rect 3476 149376 3482 149388
rect 85960 149376 85988 149484
rect 86402 149404 86408 149456
rect 86460 149404 86466 149456
rect 86420 149376 86448 149404
rect 3476 149348 85988 149376
rect 86328 149348 86448 149376
rect 86512 149376 86540 149484
rect 86678 149472 86684 149524
rect 86736 149512 86742 149524
rect 86736 149484 92060 149512
rect 86736 149472 86742 149484
rect 89438 149404 89444 149456
rect 89496 149444 89502 149456
rect 91646 149444 91652 149456
rect 89496 149416 91652 149444
rect 89496 149404 89502 149416
rect 91646 149404 91652 149416
rect 91704 149404 91710 149456
rect 91922 149404 91928 149456
rect 91980 149404 91986 149456
rect 91940 149376 91968 149404
rect 86512 149348 91968 149376
rect 3476 149336 3482 149348
rect 86328 149172 86356 149348
rect 92032 149240 92060 149484
rect 94130 149404 94136 149456
rect 94188 149404 94194 149456
rect 94148 149308 94176 149404
rect 96586 149376 96614 149552
rect 99346 149444 99374 149620
rect 118142 149540 118148 149592
rect 118200 149580 118206 149592
rect 128078 149580 128084 149592
rect 118200 149552 128084 149580
rect 118200 149540 118206 149552
rect 128078 149540 128084 149552
rect 128136 149540 128142 149592
rect 103486 149484 122834 149512
rect 103486 149444 103514 149484
rect 122558 149444 122564 149456
rect 99346 149416 103514 149444
rect 114572 149416 122564 149444
rect 114572 149376 114600 149416
rect 122558 149404 122564 149416
rect 122616 149404 122622 149456
rect 122806 149444 122834 149484
rect 580258 149444 580264 149456
rect 122806 149416 580264 149444
rect 580258 149404 580264 149416
rect 580316 149404 580322 149456
rect 96586 149348 114600 149376
rect 580626 149308 580632 149320
rect 94148 149280 580632 149308
rect 580626 149268 580632 149280
rect 580684 149268 580690 149320
rect 580534 149240 580540 149252
rect 92032 149212 580540 149240
rect 580534 149200 580540 149212
rect 580592 149200 580598 149252
rect 580442 149172 580448 149184
rect 86328 149144 580448 149172
rect 580442 149132 580448 149144
rect 580500 149132 580506 149184
rect 128998 133832 129004 133884
rect 129056 133872 129062 133884
rect 579982 133872 579988 133884
rect 129056 133844 579988 133872
rect 129056 133832 129062 133844
rect 579982 133832 579988 133844
rect 580040 133832 580046 133884
rect 3326 126420 3332 126472
rect 3384 126460 3390 126472
rect 7558 126460 7564 126472
rect 3384 126432 7564 126460
rect 3384 126420 3390 126432
rect 7558 126420 7564 126432
rect 7616 126420 7622 126472
rect 138658 118600 138664 118652
rect 138716 118640 138722 118652
rect 580166 118640 580172 118652
rect 138716 118612 580172 118640
rect 138716 118600 138722 118612
rect 580166 118600 580172 118612
rect 580224 118600 580230 118652
rect 2774 110100 2780 110152
rect 2832 110140 2838 110152
rect 4798 110140 4804 110152
rect 2832 110112 4804 110140
rect 2832 110100 2838 110112
rect 4798 110100 4804 110112
rect 4856 110100 4862 110152
rect 81894 101464 81900 101516
rect 81952 101504 81958 101516
rect 82354 101504 82360 101516
rect 81952 101476 82360 101504
rect 81952 101464 81958 101476
rect 82354 101464 82360 101476
rect 82412 101464 82418 101516
rect 113146 100796 114554 100824
rect 113146 100688 113174 100796
rect 114526 100756 114554 100796
rect 114526 100728 115934 100756
rect 103210 100660 113174 100688
rect 103210 100484 103238 100660
rect 115906 100620 115934 100728
rect 100128 100456 103238 100484
rect 109006 100592 110414 100620
rect 115906 100592 120074 100620
rect 81802 100240 81808 100292
rect 81860 100280 81866 100292
rect 81860 100252 92842 100280
rect 81860 100240 81866 100252
rect 80882 100172 80888 100224
rect 80940 100212 80946 100224
rect 92814 100212 92842 100252
rect 80940 100184 86954 100212
rect 92814 100184 94958 100212
rect 80940 100172 80946 100184
rect 81802 100104 81808 100156
rect 81860 100144 81866 100156
rect 81860 100116 86034 100144
rect 81860 100104 81866 100116
rect 77846 100036 77852 100088
rect 77904 100076 77910 100088
rect 77904 100048 84286 100076
rect 77904 100036 77910 100048
rect 80422 99968 80428 100020
rect 80480 100008 80486 100020
rect 80480 99980 83642 100008
rect 80480 99968 80486 99980
rect 83614 99952 83642 99980
rect 84258 99952 84286 100048
rect 86006 99952 86034 100116
rect 86632 100104 86638 100156
rect 86690 100104 86696 100156
rect 86926 100144 86954 100184
rect 86926 100116 93854 100144
rect 86650 100008 86678 100104
rect 90496 100076 90502 100088
rect 90146 100048 90502 100076
rect 86650 99980 86908 100008
rect 81434 99900 81440 99952
rect 81492 99940 81498 99952
rect 82354 99940 82360 99952
rect 81492 99912 82360 99940
rect 81492 99900 81498 99912
rect 82354 99900 82360 99912
rect 82412 99900 82418 99952
rect 83504 99940 83510 99952
rect 82694 99912 83510 99940
rect 81618 99832 81624 99884
rect 81676 99872 81682 99884
rect 82584 99872 82590 99884
rect 81676 99844 82590 99872
rect 81676 99832 81682 99844
rect 82584 99832 82590 99844
rect 82642 99832 82648 99884
rect 81434 99764 81440 99816
rect 81492 99804 81498 99816
rect 81894 99804 81900 99816
rect 81492 99776 81900 99804
rect 81492 99764 81498 99776
rect 81894 99764 81900 99776
rect 81952 99764 81958 99816
rect 79778 99696 79784 99748
rect 79836 99736 79842 99748
rect 82694 99736 82722 99912
rect 83504 99900 83510 99912
rect 83562 99900 83568 99952
rect 83596 99900 83602 99952
rect 83654 99900 83660 99952
rect 84056 99900 84062 99952
rect 84114 99900 84120 99952
rect 84148 99900 84154 99952
rect 84206 99900 84212 99952
rect 84240 99900 84246 99952
rect 84298 99900 84304 99952
rect 84332 99900 84338 99952
rect 84390 99900 84396 99952
rect 85160 99940 85166 99952
rect 84810 99912 85166 99940
rect 82768 99832 82774 99884
rect 82826 99832 82832 99884
rect 83044 99832 83050 99884
rect 83102 99832 83108 99884
rect 83320 99832 83326 99884
rect 83378 99872 83384 99884
rect 83378 99844 83550 99872
rect 83378 99832 83384 99844
rect 79836 99708 82722 99736
rect 79836 99696 79842 99708
rect 82786 99668 82814 99832
rect 82906 99668 82912 99680
rect 82786 99640 82912 99668
rect 82906 99628 82912 99640
rect 82964 99628 82970 99680
rect 83062 99668 83090 99832
rect 83228 99764 83234 99816
rect 83286 99764 83292 99816
rect 83246 99736 83274 99764
rect 83246 99708 83412 99736
rect 83182 99668 83188 99680
rect 83062 99640 83188 99668
rect 83182 99628 83188 99640
rect 83240 99628 83246 99680
rect 83384 99544 83412 99708
rect 83522 99680 83550 99844
rect 83780 99764 83786 99816
rect 83838 99764 83844 99816
rect 83522 99640 83556 99680
rect 83550 99628 83556 99640
rect 83608 99628 83614 99680
rect 83642 99628 83648 99680
rect 83700 99668 83706 99680
rect 83798 99668 83826 99764
rect 83700 99640 83826 99668
rect 83700 99628 83706 99640
rect 83366 99492 83372 99544
rect 83424 99492 83430 99544
rect 83826 99492 83832 99544
rect 83884 99532 83890 99544
rect 84074 99532 84102 99900
rect 84166 99748 84194 99900
rect 84350 99872 84378 99900
rect 84350 99844 84424 99872
rect 84396 99816 84424 99844
rect 84608 99832 84614 99884
rect 84666 99832 84672 99884
rect 84700 99832 84706 99884
rect 84758 99832 84764 99884
rect 84378 99764 84384 99816
rect 84436 99764 84442 99816
rect 84166 99708 84200 99748
rect 84194 99696 84200 99708
rect 84252 99696 84258 99748
rect 84470 99668 84476 99680
rect 83884 99504 84102 99532
rect 84304 99640 84476 99668
rect 83884 99492 83890 99504
rect 84304 99396 84332 99640
rect 84470 99628 84476 99640
rect 84528 99628 84534 99680
rect 84626 99600 84654 99832
rect 84396 99572 84654 99600
rect 84396 99464 84424 99572
rect 84470 99492 84476 99544
rect 84528 99532 84534 99544
rect 84718 99532 84746 99832
rect 84528 99504 84746 99532
rect 84528 99492 84534 99504
rect 84562 99464 84568 99476
rect 84396 99436 84568 99464
rect 84562 99424 84568 99436
rect 84620 99424 84626 99476
rect 84654 99424 84660 99476
rect 84712 99464 84718 99476
rect 84810 99464 84838 99912
rect 85160 99900 85166 99912
rect 85218 99900 85224 99952
rect 85988 99900 85994 99952
rect 86046 99900 86052 99952
rect 86172 99900 86178 99952
rect 86230 99900 86236 99952
rect 86264 99900 86270 99952
rect 86322 99900 86328 99952
rect 85804 99832 85810 99884
rect 85862 99832 85868 99884
rect 85896 99832 85902 99884
rect 85954 99832 85960 99884
rect 85344 99764 85350 99816
rect 85402 99764 85408 99816
rect 85620 99764 85626 99816
rect 85678 99764 85684 99816
rect 85362 99736 85390 99764
rect 85362 99708 85436 99736
rect 85408 99680 85436 99708
rect 85638 99680 85666 99764
rect 85390 99628 85396 99680
rect 85448 99628 85454 99680
rect 85638 99640 85672 99680
rect 85666 99628 85672 99640
rect 85724 99628 85730 99680
rect 85298 99560 85304 99612
rect 85356 99600 85362 99612
rect 85822 99600 85850 99832
rect 85914 99668 85942 99832
rect 86034 99668 86040 99680
rect 85914 99640 86040 99668
rect 86034 99628 86040 99640
rect 86092 99628 86098 99680
rect 85356 99572 85850 99600
rect 85356 99560 85362 99572
rect 84712 99436 84838 99464
rect 84712 99424 84718 99436
rect 84930 99424 84936 99476
rect 84988 99464 84994 99476
rect 85206 99464 85212 99476
rect 84988 99436 85212 99464
rect 84988 99424 84994 99436
rect 85206 99424 85212 99436
rect 85264 99424 85270 99476
rect 86190 99408 86218 99900
rect 86282 99816 86310 99900
rect 86586 99832 86592 99884
rect 86644 99832 86650 99884
rect 86282 99776 86316 99816
rect 86310 99764 86316 99776
rect 86368 99764 86374 99816
rect 86448 99764 86454 99816
rect 86506 99764 86512 99816
rect 86466 99612 86494 99764
rect 86604 99748 86632 99832
rect 86724 99764 86730 99816
rect 86782 99804 86788 99816
rect 86782 99764 86816 99804
rect 86586 99696 86592 99748
rect 86644 99696 86650 99748
rect 86788 99680 86816 99764
rect 86770 99628 86776 99680
rect 86828 99628 86834 99680
rect 86402 99560 86408 99612
rect 86460 99572 86494 99612
rect 86460 99560 86466 99572
rect 86678 99424 86684 99476
rect 86736 99464 86742 99476
rect 86880 99464 86908 99980
rect 87000 99900 87006 99952
rect 87058 99900 87064 99952
rect 87828 99900 87834 99952
rect 87886 99900 87892 99952
rect 88012 99900 88018 99952
rect 88070 99900 88076 99952
rect 88472 99900 88478 99952
rect 88530 99900 88536 99952
rect 88564 99900 88570 99952
rect 88622 99940 88628 99952
rect 88622 99912 88886 99940
rect 88622 99900 88628 99912
rect 87018 99532 87046 99900
rect 87552 99832 87558 99884
rect 87610 99832 87616 99884
rect 87184 99764 87190 99816
rect 87242 99764 87248 99816
rect 87276 99764 87282 99816
rect 87334 99764 87340 99816
rect 87570 99804 87598 99832
rect 87524 99776 87598 99804
rect 87202 99612 87230 99764
rect 87138 99560 87144 99612
rect 87196 99572 87230 99612
rect 87294 99600 87322 99764
rect 87524 99748 87552 99776
rect 87506 99696 87512 99748
rect 87564 99696 87570 99748
rect 87846 99680 87874 99900
rect 87846 99640 87880 99680
rect 87874 99628 87880 99640
rect 87932 99628 87938 99680
rect 87294 99572 87644 99600
rect 87196 99560 87202 99572
rect 87616 99544 87644 99572
rect 87782 99560 87788 99612
rect 87840 99560 87846 99612
rect 87414 99532 87420 99544
rect 87018 99504 87420 99532
rect 87414 99492 87420 99504
rect 87472 99492 87478 99544
rect 87598 99492 87604 99544
rect 87656 99492 87662 99544
rect 86736 99436 86908 99464
rect 86736 99424 86742 99436
rect 84838 99396 84844 99408
rect 84304 99368 84844 99396
rect 84838 99356 84844 99368
rect 84896 99356 84902 99408
rect 86190 99368 86224 99408
rect 86218 99356 86224 99368
rect 86276 99356 86282 99408
rect 87046 99288 87052 99340
rect 87104 99328 87110 99340
rect 87800 99328 87828 99560
rect 87874 99492 87880 99544
rect 87932 99532 87938 99544
rect 88030 99532 88058 99900
rect 88288 99832 88294 99884
rect 88346 99832 88352 99884
rect 88306 99680 88334 99832
rect 88490 99804 88518 99900
rect 88748 99872 88754 99884
rect 88674 99844 88754 99872
rect 88490 99776 88610 99804
rect 88306 99640 88340 99680
rect 88334 99628 88340 99640
rect 88392 99628 88398 99680
rect 88150 99560 88156 99612
rect 88208 99560 88214 99612
rect 87932 99504 88058 99532
rect 87932 99492 87938 99504
rect 88168 99396 88196 99560
rect 88426 99424 88432 99476
rect 88484 99464 88490 99476
rect 88582 99464 88610 99776
rect 88484 99436 88610 99464
rect 88674 99476 88702 99844
rect 88748 99832 88754 99844
rect 88806 99832 88812 99884
rect 88858 99600 88886 99912
rect 88932 99900 88938 99952
rect 88990 99940 88996 99952
rect 88990 99900 89024 99940
rect 89208 99900 89214 99952
rect 89266 99900 89272 99952
rect 89300 99900 89306 99952
rect 89358 99900 89364 99952
rect 89576 99900 89582 99952
rect 89634 99900 89640 99952
rect 88996 99680 89024 99900
rect 89226 99748 89254 99900
rect 89162 99696 89168 99748
rect 89220 99708 89254 99748
rect 89220 99696 89226 99708
rect 88978 99628 88984 99680
rect 89036 99628 89042 99680
rect 89318 99600 89346 99900
rect 89484 99764 89490 99816
rect 89542 99764 89548 99816
rect 89502 99736 89530 99764
rect 89456 99708 89530 99736
rect 89456 99680 89484 99708
rect 89594 99680 89622 99900
rect 89438 99628 89444 99680
rect 89496 99628 89502 99680
rect 89530 99628 89536 99680
rect 89588 99640 89622 99680
rect 89588 99628 89594 99640
rect 88858 99572 89116 99600
rect 89318 99572 89944 99600
rect 89088 99544 89116 99572
rect 89916 99544 89944 99572
rect 89070 99492 89076 99544
rect 89128 99492 89134 99544
rect 89898 99492 89904 99544
rect 89956 99492 89962 99544
rect 88674 99436 88708 99476
rect 88484 99424 88490 99436
rect 88702 99424 88708 99436
rect 88760 99424 88766 99476
rect 89346 99396 89352 99408
rect 88168 99368 89352 99396
rect 89346 99356 89352 99368
rect 89404 99356 89410 99408
rect 90146 99396 90174 100048
rect 90496 100036 90502 100048
rect 90554 100036 90560 100088
rect 93716 100036 93722 100088
rect 93774 100036 93780 100088
rect 93826 100076 93854 100116
rect 93826 100048 94682 100076
rect 91020 99980 92750 100008
rect 90312 99900 90318 99952
rect 90370 99900 90376 99952
rect 90404 99900 90410 99952
rect 90462 99900 90468 99952
rect 90588 99900 90594 99952
rect 90646 99940 90652 99952
rect 90646 99900 90680 99940
rect 90220 99832 90226 99884
rect 90278 99832 90284 99884
rect 90238 99464 90266 99832
rect 90330 99748 90358 99900
rect 90422 99872 90450 99900
rect 90422 99844 90588 99872
rect 90330 99708 90364 99748
rect 90358 99696 90364 99708
rect 90416 99696 90422 99748
rect 90560 99680 90588 99844
rect 90652 99816 90680 99900
rect 90634 99764 90640 99816
rect 90692 99764 90698 99816
rect 90542 99628 90548 99680
rect 90600 99628 90606 99680
rect 91020 99612 91048 99980
rect 92722 99952 92750 99980
rect 91232 99900 91238 99952
rect 91290 99900 91296 99952
rect 91784 99940 91790 99952
rect 91434 99912 91790 99940
rect 91250 99736 91278 99900
rect 91324 99764 91330 99816
rect 91382 99764 91388 99816
rect 91112 99708 91278 99736
rect 91002 99560 91008 99612
rect 91060 99560 91066 99612
rect 91112 99600 91140 99708
rect 91186 99628 91192 99680
rect 91244 99668 91250 99680
rect 91342 99668 91370 99764
rect 91244 99640 91370 99668
rect 91244 99628 91250 99640
rect 91278 99600 91284 99612
rect 91112 99572 91284 99600
rect 91278 99560 91284 99572
rect 91336 99560 91342 99612
rect 90726 99464 90732 99476
rect 90238 99436 90732 99464
rect 90726 99424 90732 99436
rect 90784 99424 90790 99476
rect 90818 99396 90824 99408
rect 90146 99368 90824 99396
rect 90818 99356 90824 99368
rect 90876 99356 90882 99408
rect 87104 99300 87828 99328
rect 91434 99328 91462 99912
rect 91784 99900 91790 99912
rect 91842 99900 91848 99952
rect 92336 99900 92342 99952
rect 92394 99900 92400 99952
rect 92704 99900 92710 99952
rect 92762 99900 92768 99952
rect 92888 99900 92894 99952
rect 92946 99900 92952 99952
rect 92980 99900 92986 99952
rect 93038 99900 93044 99952
rect 93256 99900 93262 99952
rect 93314 99900 93320 99952
rect 93348 99900 93354 99952
rect 93406 99900 93412 99952
rect 91508 99832 91514 99884
rect 91566 99832 91572 99884
rect 91600 99832 91606 99884
rect 91658 99832 91664 99884
rect 92152 99832 92158 99884
rect 92210 99832 92216 99884
rect 91526 99532 91554 99832
rect 91618 99612 91646 99832
rect 91618 99572 91652 99612
rect 91646 99560 91652 99572
rect 91704 99560 91710 99612
rect 92014 99560 92020 99612
rect 92072 99600 92078 99612
rect 92170 99600 92198 99832
rect 92354 99680 92382 99900
rect 92428 99832 92434 99884
rect 92486 99872 92492 99884
rect 92486 99832 92520 99872
rect 92290 99628 92296 99680
rect 92348 99640 92382 99680
rect 92348 99628 92354 99640
rect 92492 99612 92520 99832
rect 92906 99748 92934 99900
rect 92842 99696 92848 99748
rect 92900 99708 92934 99748
rect 92900 99696 92906 99708
rect 92998 99668 93026 99900
rect 93274 99872 93302 99900
rect 93228 99844 93302 99872
rect 92998 99640 93164 99668
rect 93136 99612 93164 99640
rect 93228 99612 93256 99844
rect 93366 99816 93394 99900
rect 93302 99764 93308 99816
rect 93360 99776 93394 99816
rect 93360 99764 93366 99776
rect 93394 99628 93400 99680
rect 93452 99668 93458 99680
rect 93734 99668 93762 100036
rect 93900 99900 93906 99952
rect 93958 99900 93964 99952
rect 93992 99900 93998 99952
rect 94050 99900 94056 99952
rect 93918 99680 93946 99900
rect 93452 99640 93762 99668
rect 93452 99628 93458 99640
rect 93854 99628 93860 99680
rect 93912 99640 93946 99680
rect 93912 99628 93918 99640
rect 94010 99612 94038 99900
rect 92072 99572 92198 99600
rect 92072 99560 92078 99572
rect 92474 99560 92480 99612
rect 92532 99560 92538 99612
rect 93118 99560 93124 99612
rect 93176 99560 93182 99612
rect 93210 99560 93216 99612
rect 93268 99560 93274 99612
rect 93946 99560 93952 99612
rect 94004 99572 94038 99612
rect 94004 99560 94010 99572
rect 94102 99544 94130 100048
rect 94654 99952 94682 100048
rect 94930 99952 94958 100184
rect 97580 100172 97586 100224
rect 97638 100172 97644 100224
rect 94360 99900 94366 99952
rect 94418 99900 94424 99952
rect 94636 99900 94642 99952
rect 94694 99900 94700 99952
rect 94728 99900 94734 99952
rect 94786 99900 94792 99952
rect 94912 99900 94918 99952
rect 94970 99900 94976 99952
rect 95740 99900 95746 99952
rect 95798 99900 95804 99952
rect 95924 99900 95930 99952
rect 95982 99900 95988 99952
rect 96016 99900 96022 99952
rect 96074 99900 96080 99952
rect 96292 99900 96298 99952
rect 96350 99900 96356 99952
rect 96568 99900 96574 99952
rect 96626 99940 96632 99952
rect 96626 99912 96752 99940
rect 96626 99900 96632 99912
rect 92290 99532 92296 99544
rect 91526 99504 92296 99532
rect 92290 99492 92296 99504
rect 92348 99492 92354 99544
rect 94038 99492 94044 99544
rect 94096 99504 94130 99544
rect 94096 99492 94102 99504
rect 94222 99492 94228 99544
rect 94280 99532 94286 99544
rect 94378 99532 94406 99900
rect 94544 99832 94550 99884
rect 94602 99832 94608 99884
rect 94562 99736 94590 99832
rect 94746 99816 94774 99900
rect 94682 99764 94688 99816
rect 94740 99776 94774 99816
rect 94930 99804 94958 99900
rect 95096 99832 95102 99884
rect 95154 99872 95160 99884
rect 95154 99844 95648 99872
rect 95154 99832 95160 99844
rect 94930 99776 95004 99804
rect 94740 99764 94746 99776
rect 94866 99736 94872 99748
rect 94562 99708 94872 99736
rect 94866 99696 94872 99708
rect 94924 99696 94930 99748
rect 94976 99680 95004 99776
rect 95188 99764 95194 99816
rect 95246 99764 95252 99816
rect 94958 99628 94964 99680
rect 95016 99628 95022 99680
rect 95206 99532 95234 99764
rect 94280 99504 94406 99532
rect 95068 99504 95234 99532
rect 94280 99492 94286 99504
rect 95068 99476 95096 99504
rect 93302 99424 93308 99476
rect 93360 99464 93366 99476
rect 93578 99464 93584 99476
rect 93360 99436 93584 99464
rect 93360 99424 93366 99436
rect 93578 99424 93584 99436
rect 93636 99424 93642 99476
rect 95050 99424 95056 99476
rect 95108 99424 95114 99476
rect 95142 99424 95148 99476
rect 95200 99464 95206 99476
rect 95620 99464 95648 99844
rect 95200 99436 95648 99464
rect 95200 99424 95206 99436
rect 93578 99328 93584 99340
rect 91434 99300 93584 99328
rect 87104 99288 87110 99300
rect 93578 99288 93584 99300
rect 93636 99288 93642 99340
rect 81710 99220 81716 99272
rect 81768 99260 81774 99272
rect 95758 99260 95786 99900
rect 95942 99872 95970 99900
rect 95896 99844 95970 99872
rect 95896 99680 95924 99844
rect 96034 99816 96062 99900
rect 95970 99764 95976 99816
rect 96028 99776 96062 99816
rect 96028 99764 96034 99776
rect 95878 99628 95884 99680
rect 95936 99628 95942 99680
rect 96310 99532 96338 99900
rect 96724 99680 96752 99912
rect 96936 99900 96942 99952
rect 96994 99900 97000 99952
rect 96844 99872 96850 99884
rect 96816 99832 96850 99872
rect 96902 99832 96908 99884
rect 96706 99628 96712 99680
rect 96764 99628 96770 99680
rect 96816 99668 96844 99832
rect 96954 99748 96982 99900
rect 97120 99872 97126 99884
rect 97092 99832 97126 99872
rect 97178 99832 97184 99884
rect 97304 99832 97310 99884
rect 97362 99832 97368 99884
rect 97092 99748 97120 99832
rect 96890 99696 96896 99748
rect 96948 99708 96982 99748
rect 96948 99696 96954 99708
rect 97074 99696 97080 99748
rect 97132 99696 97138 99748
rect 97166 99668 97172 99680
rect 96816 99640 97172 99668
rect 97166 99628 97172 99640
rect 97224 99628 97230 99680
rect 97322 99600 97350 99832
rect 97598 99680 97626 100172
rect 98960 100144 98966 100156
rect 98610 100116 98966 100144
rect 97672 99900 97678 99952
rect 97730 99940 97736 99952
rect 97730 99912 97902 99940
rect 97730 99900 97736 99912
rect 97764 99832 97770 99884
rect 97822 99832 97828 99884
rect 97598 99640 97632 99680
rect 97626 99628 97632 99640
rect 97684 99628 97690 99680
rect 97442 99600 97448 99612
rect 97322 99572 97448 99600
rect 97442 99560 97448 99572
rect 97500 99560 97506 99612
rect 97534 99560 97540 99612
rect 97592 99600 97598 99612
rect 97782 99600 97810 99832
rect 97592 99572 97810 99600
rect 97592 99560 97598 99572
rect 97874 99544 97902 99912
rect 97948 99900 97954 99952
rect 98006 99900 98012 99952
rect 98224 99900 98230 99952
rect 98282 99900 98288 99952
rect 98408 99940 98414 99952
rect 98380 99900 98414 99940
rect 98466 99900 98472 99952
rect 97966 99612 97994 99900
rect 98132 99764 98138 99816
rect 98190 99764 98196 99816
rect 97966 99572 98000 99612
rect 97994 99560 98000 99572
rect 98052 99560 98058 99612
rect 96430 99532 96436 99544
rect 96310 99504 96436 99532
rect 96430 99492 96436 99504
rect 96488 99492 96494 99544
rect 97874 99504 97908 99544
rect 97902 99492 97908 99504
rect 97960 99492 97966 99544
rect 98150 99396 98178 99764
rect 98242 99668 98270 99900
rect 98380 99748 98408 99900
rect 98362 99696 98368 99748
rect 98420 99696 98426 99748
rect 98454 99668 98460 99680
rect 98242 99640 98460 99668
rect 98454 99628 98460 99640
rect 98512 99628 98518 99680
rect 98610 99464 98638 100116
rect 98960 100104 98966 100116
rect 99018 100104 99024 100156
rect 100128 100144 100156 100456
rect 109006 100212 109034 100592
rect 110386 100552 110414 100592
rect 110386 100524 115934 100552
rect 99990 100116 100156 100144
rect 100358 100184 109034 100212
rect 115906 100212 115934 100524
rect 120046 100484 120074 100592
rect 120046 100456 122834 100484
rect 122806 100348 122834 100456
rect 128170 100348 128176 100360
rect 122806 100320 128176 100348
rect 128170 100308 128176 100320
rect 128228 100308 128234 100360
rect 118666 100252 120074 100280
rect 118666 100212 118694 100252
rect 115906 100184 118694 100212
rect 120046 100212 120074 100252
rect 120046 100184 125594 100212
rect 99604 100036 99610 100088
rect 99662 100076 99668 100088
rect 99662 100048 99834 100076
rect 99662 100036 99668 100048
rect 99024 99980 99696 100008
rect 98684 99900 98690 99952
rect 98742 99900 98748 99952
rect 98868 99900 98874 99952
rect 98926 99900 98932 99952
rect 98702 99748 98730 99900
rect 98886 99748 98914 99900
rect 99024 99884 99052 99980
rect 99144 99940 99150 99952
rect 99116 99900 99150 99940
rect 99202 99900 99208 99952
rect 99512 99900 99518 99952
rect 99570 99900 99576 99952
rect 99006 99832 99012 99884
rect 99064 99832 99070 99884
rect 99116 99816 99144 99900
rect 99236 99832 99242 99884
rect 99294 99832 99300 99884
rect 99420 99832 99426 99884
rect 99478 99832 99484 99884
rect 99098 99764 99104 99816
rect 99156 99764 99162 99816
rect 98702 99708 98736 99748
rect 98730 99696 98736 99708
rect 98788 99696 98794 99748
rect 98886 99708 98920 99748
rect 98914 99696 98920 99708
rect 98972 99696 98978 99748
rect 98822 99560 98828 99612
rect 98880 99600 98886 99612
rect 99254 99600 99282 99832
rect 99438 99668 99466 99832
rect 99530 99748 99558 99900
rect 99668 99816 99696 99980
rect 99650 99764 99656 99816
rect 99708 99764 99714 99816
rect 99530 99708 99564 99748
rect 99558 99696 99564 99708
rect 99616 99696 99622 99748
rect 99438 99640 99696 99668
rect 98880 99572 99282 99600
rect 98880 99560 98886 99572
rect 99006 99464 99012 99476
rect 98610 99436 99012 99464
rect 99006 99424 99012 99436
rect 99064 99424 99070 99476
rect 99668 99464 99696 99640
rect 99806 99600 99834 100048
rect 99990 99940 100018 100116
rect 100156 99940 100162 99952
rect 99990 99912 100162 99940
rect 100156 99900 100162 99912
rect 100214 99900 100220 99952
rect 100248 99900 100254 99952
rect 100306 99900 100312 99952
rect 100064 99832 100070 99884
rect 100122 99832 100128 99884
rect 100082 99736 100110 99832
rect 100266 99804 100294 99900
rect 100220 99776 100294 99804
rect 100082 99708 100156 99736
rect 99926 99600 99932 99612
rect 99806 99572 99932 99600
rect 99926 99560 99932 99572
rect 99984 99560 99990 99612
rect 99742 99492 99748 99544
rect 99800 99532 99806 99544
rect 100128 99532 100156 99708
rect 100220 99612 100248 99776
rect 100202 99560 100208 99612
rect 100260 99560 100266 99612
rect 99800 99504 100156 99532
rect 99800 99492 99806 99504
rect 99834 99464 99840 99476
rect 99668 99436 99840 99464
rect 99834 99424 99840 99436
rect 99892 99424 99898 99476
rect 100018 99424 100024 99476
rect 100076 99464 100082 99476
rect 100358 99464 100386 100184
rect 100450 100116 112714 100144
rect 100450 99952 100478 100116
rect 100708 100036 100714 100088
rect 100766 100036 100772 100088
rect 104848 100036 104854 100088
rect 104906 100036 104912 100088
rect 107332 100036 107338 100088
rect 107390 100036 107396 100088
rect 112576 100036 112582 100088
rect 112634 100036 112640 100088
rect 100726 100008 100754 100036
rect 100726 99980 101996 100008
rect 100432 99900 100438 99952
rect 100490 99900 100496 99952
rect 100616 99900 100622 99952
rect 100674 99900 100680 99952
rect 100892 99900 100898 99952
rect 100950 99900 100956 99952
rect 101076 99900 101082 99952
rect 101134 99900 101140 99952
rect 101260 99900 101266 99952
rect 101318 99900 101324 99952
rect 101444 99900 101450 99952
rect 101502 99900 101508 99952
rect 101720 99900 101726 99952
rect 101778 99940 101784 99952
rect 101778 99912 101904 99940
rect 101778 99900 101784 99912
rect 100450 99804 100478 99900
rect 100634 99816 100662 99900
rect 100450 99776 100524 99804
rect 100634 99776 100668 99816
rect 100496 99612 100524 99776
rect 100662 99764 100668 99776
rect 100720 99764 100726 99816
rect 100910 99680 100938 99900
rect 101094 99680 101122 99900
rect 100910 99640 100944 99680
rect 100938 99628 100944 99640
rect 100996 99628 101002 99680
rect 101094 99640 101128 99680
rect 101122 99628 101128 99640
rect 101180 99628 101186 99680
rect 101278 99612 101306 99900
rect 101462 99872 101490 99900
rect 101462 99844 101812 99872
rect 101536 99764 101542 99816
rect 101594 99804 101600 99816
rect 101594 99776 101720 99804
rect 101594 99764 101600 99776
rect 101582 99668 101588 99680
rect 101416 99640 101588 99668
rect 101416 99612 101444 99640
rect 101582 99628 101588 99640
rect 101640 99628 101646 99680
rect 100478 99560 100484 99612
rect 100536 99560 100542 99612
rect 101278 99572 101312 99612
rect 101306 99560 101312 99572
rect 101364 99560 101370 99612
rect 101398 99560 101404 99612
rect 101456 99560 101462 99612
rect 101490 99560 101496 99612
rect 101548 99600 101554 99612
rect 101692 99600 101720 99776
rect 101548 99572 101720 99600
rect 101548 99560 101554 99572
rect 100754 99492 100760 99544
rect 100812 99532 100818 99544
rect 101784 99532 101812 99844
rect 101876 99612 101904 99912
rect 101858 99560 101864 99612
rect 101916 99560 101922 99612
rect 101968 99544 101996 99980
rect 104038 99980 104250 100008
rect 104038 99952 104066 99980
rect 102088 99940 102094 99952
rect 102060 99900 102094 99940
rect 102146 99900 102152 99952
rect 102180 99900 102186 99952
rect 102238 99900 102244 99952
rect 102272 99900 102278 99952
rect 102330 99900 102336 99952
rect 102364 99900 102370 99952
rect 102422 99900 102428 99952
rect 102456 99900 102462 99952
rect 102514 99940 102520 99952
rect 102514 99900 102548 99940
rect 102824 99900 102830 99952
rect 102882 99940 102888 99952
rect 102882 99912 103192 99940
rect 102882 99900 102888 99912
rect 102060 99816 102088 99900
rect 102042 99764 102048 99816
rect 102100 99764 102106 99816
rect 100812 99504 101812 99532
rect 100812 99492 100818 99504
rect 101950 99492 101956 99544
rect 102008 99492 102014 99544
rect 100076 99436 100386 99464
rect 100076 99424 100082 99436
rect 101030 99396 101036 99408
rect 98150 99368 101036 99396
rect 101030 99356 101036 99368
rect 101088 99356 101094 99408
rect 102198 99396 102226 99900
rect 102290 99816 102318 99900
rect 102382 99872 102410 99900
rect 102382 99844 102456 99872
rect 102290 99776 102324 99816
rect 102318 99764 102324 99776
rect 102376 99764 102382 99816
rect 102428 99748 102456 99844
rect 102410 99696 102416 99748
rect 102468 99696 102474 99748
rect 102520 99532 102548 99900
rect 102640 99872 102646 99884
rect 102612 99832 102646 99872
rect 102698 99832 102704 99884
rect 102612 99612 102640 99832
rect 103008 99764 103014 99816
rect 103066 99764 103072 99816
rect 103026 99680 103054 99764
rect 102962 99628 102968 99680
rect 103020 99640 103054 99680
rect 103020 99628 103026 99640
rect 102594 99560 102600 99612
rect 102652 99560 102658 99612
rect 102686 99532 102692 99544
rect 102520 99504 102692 99532
rect 102686 99492 102692 99504
rect 102744 99492 102750 99544
rect 103164 99532 103192 99912
rect 103284 99900 103290 99952
rect 103342 99900 103348 99952
rect 103468 99900 103474 99952
rect 103526 99900 103532 99952
rect 103744 99900 103750 99952
rect 103802 99900 103808 99952
rect 103836 99900 103842 99952
rect 103894 99900 103900 99952
rect 103928 99900 103934 99952
rect 103986 99900 103992 99952
rect 104020 99900 104026 99952
rect 104078 99900 104084 99952
rect 104112 99900 104118 99952
rect 104170 99900 104176 99952
rect 103302 99816 103330 99900
rect 103284 99764 103290 99816
rect 103342 99764 103348 99816
rect 103376 99764 103382 99816
rect 103434 99764 103440 99816
rect 103394 99680 103422 99764
rect 103330 99628 103336 99680
rect 103388 99640 103422 99680
rect 103388 99628 103394 99640
rect 103486 99612 103514 99900
rect 103652 99832 103658 99884
rect 103710 99832 103716 99884
rect 103422 99560 103428 99612
rect 103480 99572 103514 99612
rect 103670 99600 103698 99832
rect 103624 99572 103698 99600
rect 103480 99560 103486 99572
rect 103624 99544 103652 99572
rect 103762 99544 103790 99900
rect 103854 99748 103882 99900
rect 103946 99872 103974 99900
rect 103946 99844 104020 99872
rect 103854 99708 103888 99748
rect 103882 99696 103888 99708
rect 103940 99696 103946 99748
rect 103992 99680 104020 99844
rect 104130 99680 104158 99900
rect 103974 99628 103980 99680
rect 104032 99628 104038 99680
rect 104066 99628 104072 99680
rect 104124 99640 104158 99680
rect 104124 99628 104130 99640
rect 103330 99532 103336 99544
rect 103164 99504 103336 99532
rect 103330 99492 103336 99504
rect 103388 99492 103394 99544
rect 103606 99492 103612 99544
rect 103664 99492 103670 99544
rect 103698 99492 103704 99544
rect 103756 99504 103790 99544
rect 103756 99492 103762 99504
rect 103790 99424 103796 99476
rect 103848 99464 103854 99476
rect 104222 99464 104250 99980
rect 103848 99436 104250 99464
rect 104314 99980 104710 100008
rect 103848 99424 103854 99436
rect 104314 99408 104342 99980
rect 104682 99952 104710 99980
rect 104388 99900 104394 99952
rect 104446 99900 104452 99952
rect 104664 99900 104670 99952
rect 104722 99900 104728 99952
rect 104866 99940 104894 100036
rect 104866 99912 104940 99940
rect 104406 99680 104434 99900
rect 104480 99832 104486 99884
rect 104538 99872 104544 99884
rect 104802 99872 104808 99884
rect 104538 99844 104664 99872
rect 104538 99832 104544 99844
rect 104636 99816 104664 99844
rect 104728 99844 104808 99872
rect 104618 99764 104624 99816
rect 104676 99764 104682 99816
rect 104728 99748 104756 99844
rect 104802 99832 104808 99844
rect 104860 99832 104866 99884
rect 104912 99748 104940 99912
rect 105124 99900 105130 99952
rect 105182 99900 105188 99952
rect 105308 99900 105314 99952
rect 105366 99900 105372 99952
rect 105492 99900 105498 99952
rect 105550 99900 105556 99952
rect 106228 99900 106234 99952
rect 106286 99900 106292 99952
rect 106320 99900 106326 99952
rect 106378 99900 106384 99952
rect 106504 99900 106510 99952
rect 106562 99900 106568 99952
rect 106688 99900 106694 99952
rect 106746 99900 106752 99952
rect 106872 99940 106878 99952
rect 106798 99912 106878 99940
rect 105032 99872 105038 99884
rect 105004 99832 105038 99872
rect 105090 99832 105096 99884
rect 104710 99696 104716 99748
rect 104768 99696 104774 99748
rect 104894 99696 104900 99748
rect 104952 99696 104958 99748
rect 104406 99640 104440 99680
rect 104434 99628 104440 99640
rect 104492 99628 104498 99680
rect 104802 99628 104808 99680
rect 104860 99668 104866 99680
rect 105004 99668 105032 99832
rect 104860 99640 105032 99668
rect 104860 99628 104866 99640
rect 105142 99612 105170 99900
rect 105078 99560 105084 99612
rect 105136 99572 105170 99612
rect 105136 99560 105142 99572
rect 102870 99396 102876 99408
rect 102198 99368 102876 99396
rect 102870 99356 102876 99368
rect 102928 99356 102934 99408
rect 104250 99356 104256 99408
rect 104308 99368 104342 99408
rect 105326 99396 105354 99900
rect 105400 99832 105406 99884
rect 105458 99832 105464 99884
rect 105418 99544 105446 99832
rect 105510 99680 105538 99900
rect 105952 99832 105958 99884
rect 106010 99872 106016 99884
rect 106136 99872 106142 99884
rect 106010 99832 106044 99872
rect 106016 99748 106044 99832
rect 106108 99832 106142 99872
rect 106194 99832 106200 99884
rect 105998 99696 106004 99748
rect 106056 99696 106062 99748
rect 106108 99680 106136 99832
rect 106246 99804 106274 99900
rect 106200 99776 106274 99804
rect 106200 99680 106228 99776
rect 106338 99748 106366 99900
rect 106412 99764 106418 99816
rect 106470 99764 106476 99816
rect 106274 99696 106280 99748
rect 106332 99708 106366 99748
rect 106332 99696 106338 99708
rect 105510 99640 105544 99680
rect 105538 99628 105544 99640
rect 105596 99628 105602 99680
rect 106090 99628 106096 99680
rect 106148 99628 106154 99680
rect 106182 99628 106188 99680
rect 106240 99628 106246 99680
rect 106430 99612 106458 99764
rect 106366 99560 106372 99612
rect 106424 99572 106458 99612
rect 106424 99560 106430 99572
rect 105418 99504 105452 99544
rect 105446 99492 105452 99504
rect 105504 99492 105510 99544
rect 106522 99476 106550 99900
rect 106706 99612 106734 99900
rect 106642 99560 106648 99612
rect 106700 99572 106734 99612
rect 106700 99560 106706 99572
rect 106798 99544 106826 99912
rect 106872 99900 106878 99912
rect 106930 99900 106936 99952
rect 106964 99900 106970 99952
rect 107022 99900 107028 99952
rect 107056 99900 107062 99952
rect 107114 99900 107120 99952
rect 107350 99940 107378 100036
rect 109908 100008 109914 100020
rect 109742 99980 109914 100008
rect 107350 99912 107516 99940
rect 106982 99816 107010 99900
rect 106918 99764 106924 99816
rect 106976 99776 107010 99816
rect 106976 99764 106982 99776
rect 107074 99748 107102 99900
rect 107488 99748 107516 99912
rect 107608 99900 107614 99952
rect 107666 99900 107672 99952
rect 107700 99900 107706 99952
rect 107758 99940 107764 99952
rect 107758 99900 107792 99940
rect 107976 99900 107982 99952
rect 108034 99900 108040 99952
rect 108344 99940 108350 99952
rect 108316 99900 108350 99940
rect 108402 99900 108408 99952
rect 108528 99940 108534 99952
rect 108500 99900 108534 99940
rect 108586 99900 108592 99952
rect 109080 99900 109086 99952
rect 109138 99900 109144 99952
rect 107626 99816 107654 99900
rect 107626 99776 107660 99816
rect 107654 99764 107660 99776
rect 107712 99764 107718 99816
rect 107010 99696 107016 99748
rect 107068 99708 107102 99748
rect 107068 99696 107074 99708
rect 107470 99696 107476 99748
rect 107528 99696 107534 99748
rect 107378 99560 107384 99612
rect 107436 99600 107442 99612
rect 107764 99600 107792 99900
rect 107436 99572 107792 99600
rect 107994 99600 108022 99900
rect 108114 99600 108120 99612
rect 107994 99572 108120 99600
rect 107436 99560 107442 99572
rect 108114 99560 108120 99572
rect 108172 99560 108178 99612
rect 106734 99492 106740 99544
rect 106792 99504 106826 99544
rect 108316 99532 108344 99900
rect 108390 99532 108396 99544
rect 108316 99504 108396 99532
rect 106792 99492 106798 99504
rect 108390 99492 108396 99504
rect 108448 99492 108454 99544
rect 108500 99476 108528 99900
rect 108988 99804 108994 99816
rect 108960 99764 108994 99804
rect 109046 99764 109052 99816
rect 108804 99696 108810 99748
rect 108862 99696 108868 99748
rect 108822 99600 108850 99696
rect 108960 99612 108988 99764
rect 109098 99680 109126 99900
rect 109356 99832 109362 99884
rect 109414 99832 109420 99884
rect 109034 99628 109040 99680
rect 109092 99640 109126 99680
rect 109092 99628 109098 99640
rect 108684 99572 108850 99600
rect 108684 99544 108712 99572
rect 108942 99560 108948 99612
rect 109000 99560 109006 99612
rect 108666 99492 108672 99544
rect 108724 99492 108730 99544
rect 106458 99424 106464 99476
rect 106516 99436 106550 99476
rect 106516 99424 106522 99436
rect 108482 99424 108488 99476
rect 108540 99424 108546 99476
rect 109374 99464 109402 99832
rect 109742 99532 109770 99980
rect 109908 99968 109914 99980
rect 109966 99968 109972 100020
rect 109816 99900 109822 99952
rect 109874 99900 109880 99952
rect 110000 99900 110006 99952
rect 110058 99900 110064 99952
rect 110092 99900 110098 99952
rect 110150 99900 110156 99952
rect 110460 99900 110466 99952
rect 110518 99940 110524 99952
rect 110518 99912 110736 99940
rect 110518 99900 110524 99912
rect 109834 99680 109862 99900
rect 110018 99872 110046 99900
rect 109972 99844 110046 99872
rect 109834 99640 109868 99680
rect 109862 99628 109868 99640
rect 109920 99628 109926 99680
rect 109972 99668 110000 99844
rect 110110 99804 110138 99900
rect 110276 99832 110282 99884
rect 110334 99832 110340 99884
rect 110368 99832 110374 99884
rect 110426 99872 110432 99884
rect 110426 99832 110460 99872
rect 110064 99776 110138 99804
rect 110064 99748 110092 99776
rect 110046 99696 110052 99748
rect 110104 99696 110110 99748
rect 110138 99696 110144 99748
rect 110196 99736 110202 99748
rect 110294 99736 110322 99832
rect 110432 99748 110460 99832
rect 110552 99764 110558 99816
rect 110610 99764 110616 99816
rect 110196 99708 110322 99736
rect 110196 99696 110202 99708
rect 110414 99696 110420 99748
rect 110472 99696 110478 99748
rect 110570 99680 110598 99764
rect 110230 99668 110236 99680
rect 109972 99640 110236 99668
rect 110230 99628 110236 99640
rect 110288 99628 110294 99680
rect 110506 99628 110512 99680
rect 110564 99640 110598 99680
rect 110564 99628 110570 99640
rect 110708 99544 110736 99912
rect 110828 99900 110834 99952
rect 110886 99900 110892 99952
rect 111012 99900 111018 99952
rect 111070 99900 111076 99952
rect 111104 99900 111110 99952
rect 111162 99900 111168 99952
rect 111564 99900 111570 99952
rect 111622 99940 111628 99952
rect 111622 99912 111794 99940
rect 111622 99900 111628 99912
rect 110846 99600 110874 99900
rect 111030 99668 111058 99900
rect 111122 99816 111150 99900
rect 111472 99832 111478 99884
rect 111530 99832 111536 99884
rect 111656 99832 111662 99884
rect 111714 99832 111720 99884
rect 111122 99776 111156 99816
rect 111150 99764 111156 99776
rect 111208 99764 111214 99816
rect 111490 99748 111518 99832
rect 111426 99696 111432 99748
rect 111484 99708 111518 99748
rect 111484 99696 111490 99708
rect 111674 99680 111702 99832
rect 111030 99640 111196 99668
rect 111058 99600 111064 99612
rect 110846 99572 111064 99600
rect 111058 99560 111064 99572
rect 111116 99560 111122 99612
rect 109954 99532 109960 99544
rect 109742 99504 109960 99532
rect 109954 99492 109960 99504
rect 110012 99492 110018 99544
rect 110690 99492 110696 99544
rect 110748 99492 110754 99544
rect 110874 99492 110880 99544
rect 110932 99532 110938 99544
rect 111168 99532 111196 99640
rect 111610 99628 111616 99680
rect 111668 99640 111702 99680
rect 111668 99628 111674 99640
rect 111766 99612 111794 99912
rect 112024 99900 112030 99952
rect 112082 99900 112088 99952
rect 112594 99940 112622 100036
rect 112226 99912 112622 99940
rect 111840 99832 111846 99884
rect 111898 99832 111904 99884
rect 111334 99560 111340 99612
rect 111392 99600 111398 99612
rect 111518 99600 111524 99612
rect 111392 99572 111524 99600
rect 111392 99560 111398 99572
rect 111518 99560 111524 99572
rect 111576 99560 111582 99612
rect 111702 99560 111708 99612
rect 111760 99572 111794 99612
rect 111760 99560 111766 99572
rect 110932 99504 111196 99532
rect 110932 99492 110938 99504
rect 109678 99464 109684 99476
rect 109374 99436 109684 99464
rect 109678 99424 109684 99436
rect 109736 99424 109742 99476
rect 105998 99396 106004 99408
rect 105326 99368 106004 99396
rect 104308 99356 104314 99368
rect 105998 99356 106004 99368
rect 106056 99356 106062 99408
rect 96062 99260 96068 99272
rect 81768 99232 96068 99260
rect 81768 99220 81774 99232
rect 96062 99220 96068 99232
rect 96120 99220 96126 99272
rect 111610 99220 111616 99272
rect 111668 99260 111674 99272
rect 111858 99260 111886 99832
rect 112042 99680 112070 99900
rect 111978 99628 111984 99680
rect 112036 99640 112070 99680
rect 112036 99628 112042 99640
rect 111978 99356 111984 99408
rect 112036 99396 112042 99408
rect 112226 99396 112254 99912
rect 112300 99832 112306 99884
rect 112358 99832 112364 99884
rect 112036 99368 112254 99396
rect 112318 99396 112346 99832
rect 112686 99532 112714 100116
rect 117636 100104 117642 100156
rect 117694 100104 117700 100156
rect 121592 100144 121598 100156
rect 121104 100116 121598 100144
rect 114710 100048 115842 100076
rect 113864 99968 113870 100020
rect 113922 100008 113928 100020
rect 113922 99980 114508 100008
rect 113922 99968 113928 99980
rect 113680 99940 113686 99952
rect 113422 99912 113686 99940
rect 113128 99832 113134 99884
rect 113186 99832 113192 99884
rect 113146 99600 113174 99832
rect 113266 99628 113272 99680
rect 113324 99668 113330 99680
rect 113422 99668 113450 99912
rect 113680 99900 113686 99912
rect 113738 99900 113744 99952
rect 114140 99900 114146 99952
rect 114198 99900 114204 99952
rect 113496 99832 113502 99884
rect 113554 99832 113560 99884
rect 113324 99640 113450 99668
rect 113514 99668 113542 99832
rect 114158 99736 114186 99900
rect 113836 99708 114186 99736
rect 113836 99680 113864 99708
rect 113634 99668 113640 99680
rect 113514 99640 113640 99668
rect 113324 99628 113330 99640
rect 113634 99628 113640 99640
rect 113692 99628 113698 99680
rect 113818 99628 113824 99680
rect 113876 99628 113882 99680
rect 113910 99628 113916 99680
rect 113968 99668 113974 99680
rect 114094 99668 114100 99680
rect 113968 99640 114100 99668
rect 113968 99628 113974 99640
rect 114094 99628 114100 99640
rect 114152 99628 114158 99680
rect 113450 99600 113456 99612
rect 113146 99572 113456 99600
rect 113450 99560 113456 99572
rect 113508 99560 113514 99612
rect 112686 99504 113174 99532
rect 112622 99396 112628 99408
rect 112318 99368 112628 99396
rect 112036 99356 112042 99368
rect 112622 99356 112628 99368
rect 112680 99356 112686 99408
rect 111668 99232 111886 99260
rect 113146 99260 113174 99504
rect 114480 99476 114508 99980
rect 114710 99952 114738 100048
rect 114894 99980 115290 100008
rect 114894 99952 114922 99980
rect 114692 99900 114698 99952
rect 114750 99900 114756 99952
rect 114876 99900 114882 99952
rect 114934 99900 114940 99952
rect 115152 99900 115158 99952
rect 115210 99900 115216 99952
rect 114968 99832 114974 99884
rect 115026 99832 115032 99884
rect 114986 99736 115014 99832
rect 114756 99708 115014 99736
rect 114462 99424 114468 99476
rect 114520 99424 114526 99476
rect 114756 99340 114784 99708
rect 115170 99680 115198 99900
rect 115106 99628 115112 99680
rect 115164 99640 115198 99680
rect 115164 99628 115170 99640
rect 115014 99560 115020 99612
rect 115072 99600 115078 99612
rect 115262 99600 115290 99980
rect 115336 99900 115342 99952
rect 115394 99900 115400 99952
rect 115428 99900 115434 99952
rect 115486 99900 115492 99952
rect 115072 99572 115290 99600
rect 115072 99560 115078 99572
rect 115354 99544 115382 99900
rect 115446 99680 115474 99900
rect 115704 99764 115710 99816
rect 115762 99764 115768 99816
rect 115446 99640 115480 99680
rect 115474 99628 115480 99640
rect 115532 99628 115538 99680
rect 115722 99544 115750 99764
rect 114922 99492 114928 99544
rect 114980 99532 114986 99544
rect 115198 99532 115204 99544
rect 114980 99504 115204 99532
rect 114980 99492 114986 99504
rect 115198 99492 115204 99504
rect 115256 99492 115262 99544
rect 115354 99504 115388 99544
rect 115382 99492 115388 99504
rect 115440 99492 115446 99544
rect 115658 99492 115664 99544
rect 115716 99504 115750 99544
rect 115814 99544 115842 100048
rect 116366 100048 116762 100076
rect 115888 99900 115894 99952
rect 115946 99900 115952 99952
rect 115980 99900 115986 99952
rect 116038 99900 116044 99952
rect 116072 99900 116078 99952
rect 116130 99900 116136 99952
rect 115906 99600 115934 99900
rect 115998 99668 116026 99900
rect 116090 99748 116118 99900
rect 116256 99832 116262 99884
rect 116314 99832 116320 99884
rect 116090 99708 116124 99748
rect 116118 99696 116124 99708
rect 116176 99696 116182 99748
rect 116274 99680 116302 99832
rect 116366 99736 116394 100048
rect 116734 99952 116762 100048
rect 117148 100048 117590 100076
rect 116440 99900 116446 99952
rect 116498 99900 116504 99952
rect 116624 99900 116630 99952
rect 116682 99900 116688 99952
rect 116716 99900 116722 99952
rect 116774 99900 116780 99952
rect 116808 99900 116814 99952
rect 116866 99900 116872 99952
rect 116992 99900 116998 99952
rect 117050 99940 117056 99952
rect 117050 99900 117084 99940
rect 116458 99816 116486 99900
rect 116458 99776 116492 99816
rect 116486 99764 116492 99776
rect 116544 99764 116550 99816
rect 116642 99804 116670 99900
rect 116826 99872 116854 99900
rect 116826 99844 116992 99872
rect 116642 99776 116900 99804
rect 116578 99736 116584 99748
rect 116366 99708 116584 99736
rect 116578 99696 116584 99708
rect 116636 99696 116642 99748
rect 116872 99680 116900 99776
rect 115998 99640 116164 99668
rect 116274 99640 116308 99680
rect 116026 99600 116032 99612
rect 115906 99572 116032 99600
rect 116026 99560 116032 99572
rect 116084 99560 116090 99612
rect 115814 99504 115848 99544
rect 115716 99492 115722 99504
rect 115842 99492 115848 99504
rect 115900 99492 115906 99544
rect 115934 99492 115940 99544
rect 115992 99532 115998 99544
rect 116136 99532 116164 99640
rect 116302 99628 116308 99640
rect 116360 99628 116366 99680
rect 116854 99628 116860 99680
rect 116912 99628 116918 99680
rect 116762 99560 116768 99612
rect 116820 99600 116826 99612
rect 116964 99600 116992 99844
rect 116820 99572 116992 99600
rect 116820 99560 116826 99572
rect 115992 99504 116164 99532
rect 115992 99492 115998 99504
rect 117056 99464 117084 99900
rect 117148 99680 117176 100048
rect 117562 99952 117590 100048
rect 117360 99900 117366 99952
rect 117418 99900 117424 99952
rect 117452 99900 117458 99952
rect 117510 99900 117516 99952
rect 117544 99900 117550 99952
rect 117602 99900 117608 99952
rect 117268 99832 117274 99884
rect 117326 99832 117332 99884
rect 117130 99628 117136 99680
rect 117188 99628 117194 99680
rect 117286 99532 117314 99832
rect 117378 99612 117406 99900
rect 117470 99748 117498 99900
rect 117654 99804 117682 100104
rect 117820 99940 117826 99952
rect 117608 99776 117682 99804
rect 117792 99900 117826 99940
rect 117878 99900 117884 99952
rect 117912 99900 117918 99952
rect 117970 99900 117976 99952
rect 118372 99900 118378 99952
rect 118430 99900 118436 99952
rect 118648 99900 118654 99952
rect 118706 99940 118712 99952
rect 118706 99912 119016 99940
rect 118706 99900 118712 99912
rect 117470 99708 117504 99748
rect 117498 99696 117504 99708
rect 117556 99696 117562 99748
rect 117378 99572 117412 99612
rect 117406 99560 117412 99572
rect 117464 99560 117470 99612
rect 117498 99532 117504 99544
rect 117286 99504 117504 99532
rect 117498 99492 117504 99504
rect 117556 99492 117562 99544
rect 117222 99464 117228 99476
rect 117056 99436 117228 99464
rect 117222 99424 117228 99436
rect 117280 99424 117286 99476
rect 117314 99424 117320 99476
rect 117372 99464 117378 99476
rect 117608 99464 117636 99776
rect 117682 99696 117688 99748
rect 117740 99696 117746 99748
rect 117372 99436 117636 99464
rect 117700 99464 117728 99696
rect 117792 99544 117820 99900
rect 117930 99680 117958 99900
rect 118004 99832 118010 99884
rect 118062 99832 118068 99884
rect 118188 99832 118194 99884
rect 118246 99832 118252 99884
rect 117866 99628 117872 99680
rect 117924 99640 117958 99680
rect 117924 99628 117930 99640
rect 118022 99612 118050 99832
rect 118206 99748 118234 99832
rect 118206 99708 118240 99748
rect 118234 99696 118240 99708
rect 118292 99696 118298 99748
rect 117958 99560 117964 99612
rect 118016 99572 118050 99612
rect 118390 99612 118418 99900
rect 118740 99832 118746 99884
rect 118798 99832 118804 99884
rect 118390 99572 118424 99612
rect 118016 99560 118022 99572
rect 118418 99560 118424 99572
rect 118476 99560 118482 99612
rect 118758 99544 118786 99832
rect 118988 99612 119016 99912
rect 119200 99900 119206 99952
rect 119258 99900 119264 99952
rect 119476 99900 119482 99952
rect 119534 99900 119540 99952
rect 119568 99900 119574 99952
rect 119626 99900 119632 99952
rect 119660 99900 119666 99952
rect 119718 99940 119724 99952
rect 119718 99900 119752 99940
rect 120028 99900 120034 99952
rect 120086 99900 120092 99952
rect 120120 99900 120126 99952
rect 120178 99900 120184 99952
rect 120488 99900 120494 99952
rect 120546 99900 120552 99952
rect 120580 99900 120586 99952
rect 120638 99900 120644 99952
rect 120672 99900 120678 99952
rect 120730 99900 120736 99952
rect 120948 99900 120954 99952
rect 121006 99900 121012 99952
rect 118970 99560 118976 99612
rect 119028 99560 119034 99612
rect 119218 99600 119246 99900
rect 119494 99816 119522 99900
rect 119586 99872 119614 99900
rect 119586 99844 119660 99872
rect 119632 99816 119660 99844
rect 119724 99816 119752 99900
rect 119844 99872 119850 99884
rect 119816 99832 119850 99872
rect 119902 99832 119908 99884
rect 119936 99832 119942 99884
rect 119994 99832 120000 99884
rect 119292 99764 119298 99816
rect 119350 99764 119356 99816
rect 119494 99776 119528 99816
rect 119522 99764 119528 99776
rect 119580 99764 119586 99816
rect 119614 99764 119620 99816
rect 119672 99764 119678 99816
rect 119706 99764 119712 99816
rect 119764 99764 119770 99816
rect 119310 99736 119338 99764
rect 119816 99748 119844 99832
rect 119310 99708 119660 99736
rect 119632 99680 119660 99708
rect 119798 99696 119804 99748
rect 119856 99696 119862 99748
rect 119954 99680 119982 99832
rect 119614 99628 119620 99680
rect 119672 99628 119678 99680
rect 119890 99628 119896 99680
rect 119948 99640 119982 99680
rect 119948 99628 119954 99640
rect 120046 99600 120074 99900
rect 120138 99668 120166 99900
rect 120506 99748 120534 99900
rect 120598 99804 120626 99900
rect 120690 99872 120718 99900
rect 120690 99844 120764 99872
rect 120736 99816 120764 99844
rect 120598 99776 120672 99804
rect 120644 99748 120672 99776
rect 120718 99764 120724 99816
rect 120776 99764 120782 99816
rect 120506 99708 120540 99748
rect 120534 99696 120540 99708
rect 120592 99696 120598 99748
rect 120626 99696 120632 99748
rect 120684 99696 120690 99748
rect 120810 99668 120816 99680
rect 120138 99640 120816 99668
rect 120810 99628 120816 99640
rect 120868 99628 120874 99680
rect 120166 99600 120172 99612
rect 119218 99572 119476 99600
rect 120046 99572 120172 99600
rect 117774 99492 117780 99544
rect 117832 99492 117838 99544
rect 118758 99504 118792 99544
rect 118786 99492 118792 99504
rect 118844 99492 118850 99544
rect 119448 99476 119476 99572
rect 120166 99560 120172 99572
rect 120224 99560 120230 99612
rect 120966 99476 120994 99900
rect 121104 99600 121132 100116
rect 121592 100104 121598 100116
rect 121650 100104 121656 100156
rect 125566 100144 125594 100184
rect 127986 100144 127992 100156
rect 125566 100116 127992 100144
rect 127986 100104 127992 100116
rect 128044 100104 128050 100156
rect 121316 100036 121322 100088
rect 121374 100036 121380 100088
rect 125732 100036 125738 100088
rect 125790 100036 125796 100088
rect 127112 100036 127118 100088
rect 127170 100076 127176 100088
rect 127802 100076 127808 100088
rect 127170 100048 127808 100076
rect 127170 100036 127176 100048
rect 127802 100036 127808 100048
rect 127860 100036 127866 100088
rect 121224 99764 121230 99816
rect 121282 99764 121288 99816
rect 121242 99680 121270 99764
rect 121178 99628 121184 99680
rect 121236 99640 121270 99680
rect 121334 99668 121362 100036
rect 122788 99968 122794 100020
rect 122846 99968 122852 100020
rect 124720 99968 124726 100020
rect 124778 100008 124784 100020
rect 125750 100008 125778 100036
rect 124778 99968 124812 100008
rect 125750 99980 125962 100008
rect 121408 99900 121414 99952
rect 121466 99940 121472 99952
rect 121466 99912 122144 99940
rect 121466 99900 121472 99912
rect 121868 99872 121874 99884
rect 121748 99844 121874 99872
rect 121546 99668 121552 99680
rect 121334 99640 121552 99668
rect 121236 99628 121242 99640
rect 121546 99628 121552 99640
rect 121604 99628 121610 99680
rect 121454 99600 121460 99612
rect 121104 99572 121460 99600
rect 121454 99560 121460 99572
rect 121512 99560 121518 99612
rect 121748 99544 121776 99844
rect 121868 99832 121874 99844
rect 121926 99832 121932 99884
rect 121730 99492 121736 99544
rect 121788 99492 121794 99544
rect 122116 99532 122144 99912
rect 122236 99900 122242 99952
rect 122294 99900 122300 99952
rect 122328 99900 122334 99952
rect 122386 99940 122392 99952
rect 122386 99912 122650 99940
rect 122386 99900 122392 99912
rect 122254 99668 122282 99900
rect 122374 99668 122380 99680
rect 122254 99640 122380 99668
rect 122374 99628 122380 99640
rect 122432 99628 122438 99680
rect 122282 99560 122288 99612
rect 122340 99600 122346 99612
rect 122622 99600 122650 99912
rect 122696 99900 122702 99952
rect 122754 99900 122760 99952
rect 122340 99572 122650 99600
rect 122340 99560 122346 99572
rect 122714 99544 122742 99900
rect 122116 99504 122604 99532
rect 118326 99464 118332 99476
rect 117700 99436 118332 99464
rect 117372 99424 117378 99436
rect 118326 99424 118332 99436
rect 118384 99424 118390 99476
rect 119430 99424 119436 99476
rect 119488 99424 119494 99476
rect 120966 99436 121000 99476
rect 120994 99424 121000 99436
rect 121052 99424 121058 99476
rect 122576 99464 122604 99504
rect 122650 99492 122656 99544
rect 122708 99504 122742 99544
rect 122806 99532 122834 99968
rect 123248 99900 123254 99952
rect 123306 99900 123312 99952
rect 123432 99900 123438 99952
rect 123490 99900 123496 99952
rect 123524 99900 123530 99952
rect 123582 99940 123588 99952
rect 123582 99912 123846 99940
rect 123582 99900 123588 99912
rect 123064 99832 123070 99884
rect 123122 99832 123128 99884
rect 122926 99628 122932 99680
rect 122984 99668 122990 99680
rect 123082 99668 123110 99832
rect 122984 99640 123110 99668
rect 123266 99680 123294 99900
rect 123266 99640 123300 99680
rect 122984 99628 122990 99640
rect 123294 99628 123300 99640
rect 123352 99628 123358 99680
rect 123110 99560 123116 99612
rect 123168 99600 123174 99612
rect 123450 99600 123478 99900
rect 123708 99832 123714 99884
rect 123766 99832 123772 99884
rect 123168 99572 123478 99600
rect 123168 99560 123174 99572
rect 123570 99532 123576 99544
rect 122806 99504 123576 99532
rect 122708 99492 122714 99504
rect 123570 99492 123576 99504
rect 123628 99492 123634 99544
rect 122742 99464 122748 99476
rect 122576 99436 122748 99464
rect 122742 99424 122748 99436
rect 122800 99424 122806 99476
rect 123386 99424 123392 99476
rect 123444 99464 123450 99476
rect 123726 99464 123754 99832
rect 123818 99680 123846 99912
rect 123984 99900 123990 99952
rect 124042 99900 124048 99952
rect 124076 99900 124082 99952
rect 124134 99900 124140 99952
rect 124002 99804 124030 99900
rect 123956 99776 124030 99804
rect 123956 99680 123984 99776
rect 124094 99748 124122 99900
rect 124168 99832 124174 99884
rect 124226 99832 124232 99884
rect 124352 99832 124358 99884
rect 124410 99872 124416 99884
rect 124410 99844 124720 99872
rect 124410 99832 124416 99844
rect 124030 99696 124036 99748
rect 124088 99708 124122 99748
rect 124088 99696 124094 99708
rect 123818 99640 123852 99680
rect 123846 99628 123852 99640
rect 123904 99628 123910 99680
rect 123938 99628 123944 99680
rect 123996 99628 124002 99680
rect 124186 99668 124214 99832
rect 124692 99816 124720 99844
rect 124674 99764 124680 99816
rect 124732 99764 124738 99816
rect 124306 99696 124312 99748
rect 124364 99736 124370 99748
rect 124398 99736 124404 99748
rect 124364 99708 124404 99736
rect 124364 99696 124370 99708
rect 124398 99696 124404 99708
rect 124456 99696 124462 99748
rect 124490 99668 124496 99680
rect 124186 99640 124496 99668
rect 124490 99628 124496 99640
rect 124548 99628 124554 99680
rect 124214 99492 124220 99544
rect 124272 99532 124278 99544
rect 124784 99532 124812 99968
rect 125548 99900 125554 99952
rect 125606 99900 125612 99952
rect 125566 99872 125594 99900
rect 125566 99844 125732 99872
rect 124272 99504 124812 99532
rect 124876 99708 125594 99736
rect 124272 99492 124278 99504
rect 123444 99436 123754 99464
rect 123444 99424 123450 99436
rect 124876 99396 124904 99708
rect 114848 99368 124904 99396
rect 114738 99288 114744 99340
rect 114796 99288 114802 99340
rect 114848 99260 114876 99368
rect 116486 99288 116492 99340
rect 116544 99288 116550 99340
rect 125566 99328 125594 99708
rect 125704 99408 125732 99844
rect 125824 99764 125830 99816
rect 125882 99764 125888 99816
rect 125842 99532 125870 99764
rect 125934 99612 125962 99980
rect 126946 99980 127388 100008
rect 126946 99952 126974 99980
rect 126008 99900 126014 99952
rect 126066 99900 126072 99952
rect 126284 99900 126290 99952
rect 126342 99900 126348 99952
rect 126376 99900 126382 99952
rect 126434 99900 126440 99952
rect 126928 99900 126934 99952
rect 126986 99900 126992 99952
rect 127020 99900 127026 99952
rect 127078 99900 127084 99952
rect 127204 99900 127210 99952
rect 127262 99900 127268 99952
rect 126026 99668 126054 99900
rect 126302 99748 126330 99900
rect 126394 99804 126422 99900
rect 126836 99832 126842 99884
rect 126894 99832 126900 99884
rect 126394 99776 126606 99804
rect 126238 99696 126244 99748
rect 126296 99708 126330 99748
rect 126296 99696 126302 99708
rect 126026 99640 126376 99668
rect 125934 99572 125968 99612
rect 125962 99560 125968 99572
rect 126020 99560 126026 99612
rect 126238 99532 126244 99544
rect 125842 99504 126244 99532
rect 126238 99492 126244 99504
rect 126296 99492 126302 99544
rect 126348 99532 126376 99640
rect 126422 99560 126428 99612
rect 126480 99600 126486 99612
rect 126578 99600 126606 99776
rect 126480 99572 126606 99600
rect 126854 99612 126882 99832
rect 127038 99748 127066 99900
rect 127038 99708 127072 99748
rect 127066 99696 127072 99708
rect 127124 99696 127130 99748
rect 127222 99612 127250 99900
rect 127360 99872 127388 99980
rect 127618 99872 127624 99884
rect 127360 99844 127624 99872
rect 127618 99832 127624 99844
rect 127676 99832 127682 99884
rect 126854 99572 126888 99612
rect 126480 99560 126486 99572
rect 126882 99560 126888 99572
rect 126940 99560 126946 99612
rect 127222 99572 127256 99612
rect 127250 99560 127256 99572
rect 127308 99560 127314 99612
rect 126514 99532 126520 99544
rect 126348 99504 126520 99532
rect 126514 99492 126520 99504
rect 126572 99492 126578 99544
rect 125686 99356 125692 99408
rect 125744 99356 125750 99408
rect 126146 99356 126152 99408
rect 126204 99396 126210 99408
rect 126422 99396 126428 99408
rect 126204 99368 126428 99396
rect 126204 99356 126210 99368
rect 126422 99356 126428 99368
rect 126480 99356 126486 99408
rect 128078 99328 128084 99340
rect 125566 99300 128084 99328
rect 128078 99288 128084 99300
rect 128136 99288 128142 99340
rect 113146 99232 114876 99260
rect 111668 99220 111674 99232
rect 116504 99124 116532 99288
rect 116670 99124 116676 99136
rect 116504 99096 116676 99124
rect 116670 99084 116676 99096
rect 116728 99084 116734 99136
rect 120074 98540 120080 98592
rect 120132 98580 120138 98592
rect 121362 98580 121368 98592
rect 120132 98552 121368 98580
rect 120132 98540 120138 98552
rect 121362 98540 121368 98552
rect 121420 98540 121426 98592
rect 88610 98472 88616 98524
rect 88668 98512 88674 98524
rect 88886 98512 88892 98524
rect 88668 98484 88892 98512
rect 88668 98472 88674 98484
rect 88886 98472 88892 98484
rect 88944 98472 88950 98524
rect 95234 98472 95240 98524
rect 95292 98512 95298 98524
rect 95418 98512 95424 98524
rect 95292 98484 95424 98512
rect 95292 98472 95298 98484
rect 95418 98472 95424 98484
rect 95476 98472 95482 98524
rect 89254 98336 89260 98388
rect 89312 98376 89318 98388
rect 90910 98376 90916 98388
rect 89312 98348 90916 98376
rect 89312 98336 89318 98348
rect 90910 98336 90916 98348
rect 90968 98336 90974 98388
rect 102042 98336 102048 98388
rect 102100 98376 102106 98388
rect 103238 98376 103244 98388
rect 102100 98348 103244 98376
rect 102100 98336 102106 98348
rect 103238 98336 103244 98348
rect 103296 98336 103302 98388
rect 82722 98268 82728 98320
rect 82780 98308 82786 98320
rect 86586 98308 86592 98320
rect 82780 98280 86592 98308
rect 82780 98268 82786 98280
rect 86586 98268 86592 98280
rect 86644 98268 86650 98320
rect 89714 98268 89720 98320
rect 89772 98308 89778 98320
rect 89898 98308 89904 98320
rect 89772 98280 89904 98308
rect 89772 98268 89778 98280
rect 89898 98268 89904 98280
rect 89956 98268 89962 98320
rect 117130 98268 117136 98320
rect 117188 98308 117194 98320
rect 117590 98308 117596 98320
rect 117188 98280 117596 98308
rect 117188 98268 117194 98280
rect 117590 98268 117596 98280
rect 117648 98268 117654 98320
rect 127342 98268 127348 98320
rect 127400 98308 127406 98320
rect 127710 98308 127716 98320
rect 127400 98280 127716 98308
rect 127400 98268 127406 98280
rect 127710 98268 127716 98280
rect 127768 98268 127774 98320
rect 83366 98132 83372 98184
rect 83424 98172 83430 98184
rect 83918 98172 83924 98184
rect 83424 98144 83924 98172
rect 83424 98132 83430 98144
rect 83918 98132 83924 98144
rect 83976 98132 83982 98184
rect 89438 98132 89444 98184
rect 89496 98172 89502 98184
rect 89714 98172 89720 98184
rect 89496 98144 89720 98172
rect 89496 98132 89502 98144
rect 89714 98132 89720 98144
rect 89772 98132 89778 98184
rect 91462 98132 91468 98184
rect 91520 98172 91526 98184
rect 91520 98144 92796 98172
rect 91520 98132 91526 98144
rect 90082 98064 90088 98116
rect 90140 98104 90146 98116
rect 91738 98104 91744 98116
rect 90140 98076 91744 98104
rect 90140 98064 90146 98076
rect 91738 98064 91744 98076
rect 91796 98064 91802 98116
rect 92768 97968 92796 98144
rect 103606 98132 103612 98184
rect 103664 98172 103670 98184
rect 103790 98172 103796 98184
rect 103664 98144 103796 98172
rect 103664 98132 103670 98144
rect 103790 98132 103796 98144
rect 103848 98132 103854 98184
rect 110966 98064 110972 98116
rect 111024 98104 111030 98116
rect 114278 98104 114284 98116
rect 111024 98076 114284 98104
rect 111024 98064 111030 98076
rect 114278 98064 114284 98076
rect 114336 98064 114342 98116
rect 92768 97940 109034 97968
rect 91094 97860 91100 97912
rect 91152 97900 91158 97912
rect 92106 97900 92112 97912
rect 91152 97872 92112 97900
rect 91152 97860 91158 97872
rect 92106 97860 92112 97872
rect 92164 97860 92170 97912
rect 92382 97860 92388 97912
rect 92440 97900 92446 97912
rect 109006 97900 109034 97940
rect 110966 97928 110972 97980
rect 111024 97968 111030 97980
rect 111150 97968 111156 97980
rect 111024 97940 111156 97968
rect 111024 97928 111030 97940
rect 111150 97928 111156 97940
rect 111208 97928 111214 97980
rect 113082 97928 113088 97980
rect 113140 97968 113146 97980
rect 113818 97968 113824 97980
rect 113140 97940 113824 97968
rect 113140 97928 113146 97940
rect 113818 97928 113824 97940
rect 113876 97928 113882 97980
rect 117958 97928 117964 97980
rect 118016 97968 118022 97980
rect 129182 97968 129188 97980
rect 118016 97940 129188 97968
rect 118016 97928 118022 97940
rect 129182 97928 129188 97940
rect 129240 97928 129246 97980
rect 129734 97900 129740 97912
rect 92440 97872 99374 97900
rect 109006 97872 129740 97900
rect 92440 97860 92446 97872
rect 82078 97792 82084 97844
rect 82136 97832 82142 97844
rect 82136 97804 92060 97832
rect 82136 97792 82142 97804
rect 92032 97776 92060 97804
rect 98454 97792 98460 97844
rect 98512 97832 98518 97844
rect 98822 97832 98828 97844
rect 98512 97804 98828 97832
rect 98512 97792 98518 97804
rect 98822 97792 98828 97804
rect 98880 97792 98886 97844
rect 99346 97832 99374 97872
rect 129734 97860 129740 97872
rect 129792 97860 129798 97912
rect 131114 97832 131120 97844
rect 99346 97804 131120 97832
rect 131114 97792 131120 97804
rect 131172 97792 131178 97844
rect 81986 97724 81992 97776
rect 82044 97764 82050 97776
rect 82044 97736 85574 97764
rect 82044 97724 82050 97736
rect 64874 97656 64880 97708
rect 64932 97696 64938 97708
rect 81802 97696 81808 97708
rect 64932 97668 81808 97696
rect 64932 97656 64938 97668
rect 81802 97656 81808 97668
rect 81860 97656 81866 97708
rect 62758 97588 62764 97640
rect 62816 97628 62822 97640
rect 84286 97628 84292 97640
rect 62816 97600 84292 97628
rect 62816 97588 62822 97600
rect 84286 97588 84292 97600
rect 84344 97588 84350 97640
rect 58618 97520 58624 97572
rect 58676 97560 58682 97572
rect 84378 97560 84384 97572
rect 58676 97532 84384 97560
rect 58676 97520 58682 97532
rect 84378 97520 84384 97532
rect 84436 97520 84442 97572
rect 85546 97560 85574 97736
rect 92014 97724 92020 97776
rect 92072 97764 92078 97776
rect 92382 97764 92388 97776
rect 92072 97736 92388 97764
rect 92072 97724 92078 97736
rect 92382 97724 92388 97736
rect 92440 97724 92446 97776
rect 131758 97764 131764 97776
rect 93458 97736 131764 97764
rect 89990 97656 89996 97708
rect 90048 97696 90054 97708
rect 91094 97696 91100 97708
rect 90048 97668 91100 97696
rect 90048 97656 90054 97668
rect 91094 97656 91100 97668
rect 91152 97656 91158 97708
rect 91646 97656 91652 97708
rect 91704 97696 91710 97708
rect 93458 97696 93486 97736
rect 131758 97724 131764 97736
rect 131816 97724 131822 97776
rect 91704 97668 93486 97696
rect 91704 97656 91710 97668
rect 93578 97656 93584 97708
rect 93636 97696 93642 97708
rect 133874 97696 133880 97708
rect 93636 97668 133880 97696
rect 93636 97656 93642 97668
rect 133874 97656 133880 97668
rect 133932 97656 133938 97708
rect 88426 97588 88432 97640
rect 88484 97628 88490 97640
rect 89070 97628 89076 97640
rect 88484 97600 89076 97628
rect 88484 97588 88490 97600
rect 89070 97588 89076 97600
rect 89128 97588 89134 97640
rect 92198 97588 92204 97640
rect 92256 97628 92262 97640
rect 135898 97628 135904 97640
rect 92256 97600 135904 97628
rect 92256 97588 92262 97600
rect 135898 97588 135904 97600
rect 135956 97588 135962 97640
rect 92474 97560 92480 97572
rect 85546 97532 92480 97560
rect 92474 97520 92480 97532
rect 92532 97520 92538 97572
rect 92842 97520 92848 97572
rect 92900 97560 92906 97572
rect 93486 97560 93492 97572
rect 92900 97532 93492 97560
rect 92900 97520 92906 97532
rect 93486 97520 93492 97532
rect 93544 97520 93550 97572
rect 98546 97520 98552 97572
rect 98604 97560 98610 97572
rect 99190 97560 99196 97572
rect 98604 97532 99196 97560
rect 98604 97520 98610 97532
rect 99190 97520 99196 97532
rect 99248 97520 99254 97572
rect 104894 97520 104900 97572
rect 104952 97560 104958 97572
rect 113818 97560 113824 97572
rect 104952 97532 113824 97560
rect 104952 97520 104958 97532
rect 113818 97520 113824 97532
rect 113876 97520 113882 97572
rect 118142 97560 118148 97572
rect 115906 97532 118148 97560
rect 53098 97452 53104 97504
rect 53156 97492 53162 97504
rect 79778 97492 79784 97504
rect 53156 97464 79784 97492
rect 53156 97452 53162 97464
rect 79778 97452 79784 97464
rect 79836 97452 79842 97504
rect 85758 97452 85764 97504
rect 85816 97492 85822 97504
rect 86126 97492 86132 97504
rect 85816 97464 86132 97492
rect 85816 97452 85822 97464
rect 86126 97452 86132 97464
rect 86184 97452 86190 97504
rect 106182 97452 106188 97504
rect 106240 97492 106246 97504
rect 113910 97492 113916 97504
rect 106240 97464 113916 97492
rect 106240 97452 106246 97464
rect 113910 97452 113916 97464
rect 113968 97452 113974 97504
rect 54478 97384 54484 97436
rect 54536 97424 54542 97436
rect 77846 97424 77852 97436
rect 54536 97396 77852 97424
rect 54536 97384 54542 97396
rect 77846 97384 77852 97396
rect 77904 97384 77910 97436
rect 84378 97384 84384 97436
rect 84436 97424 84442 97436
rect 86402 97424 86408 97436
rect 84436 97396 86408 97424
rect 84436 97384 84442 97396
rect 86402 97384 86408 97396
rect 86460 97384 86466 97436
rect 90818 97384 90824 97436
rect 90876 97424 90882 97436
rect 92014 97424 92020 97436
rect 90876 97396 92020 97424
rect 90876 97384 90882 97396
rect 92014 97384 92020 97396
rect 92072 97384 92078 97436
rect 101950 97384 101956 97436
rect 102008 97424 102014 97436
rect 115906 97424 115934 97532
rect 118142 97520 118148 97532
rect 118200 97520 118206 97572
rect 121362 97520 121368 97572
rect 121420 97560 121426 97572
rect 200758 97560 200764 97572
rect 121420 97532 200764 97560
rect 121420 97520 121426 97532
rect 200758 97520 200764 97532
rect 200816 97520 200822 97572
rect 127066 97452 127072 97504
rect 127124 97492 127130 97504
rect 209038 97492 209044 97504
rect 127124 97464 209044 97492
rect 127124 97452 127130 97464
rect 209038 97452 209044 97464
rect 209096 97452 209102 97504
rect 102008 97396 115934 97424
rect 102008 97384 102014 97396
rect 118970 97384 118976 97436
rect 119028 97424 119034 97436
rect 119338 97424 119344 97436
rect 119028 97396 119344 97424
rect 119028 97384 119034 97396
rect 119338 97384 119344 97396
rect 119396 97384 119402 97436
rect 122742 97384 122748 97436
rect 122800 97424 122806 97436
rect 278038 97424 278044 97436
rect 122800 97396 278044 97424
rect 122800 97384 122806 97396
rect 278038 97384 278044 97396
rect 278096 97384 278102 97436
rect 43438 97316 43444 97368
rect 43496 97356 43502 97368
rect 80422 97356 80428 97368
rect 43496 97328 80428 97356
rect 43496 97316 43502 97328
rect 80422 97316 80428 97328
rect 80480 97316 80486 97368
rect 116394 97356 116400 97368
rect 99346 97328 116400 97356
rect 31018 97248 31024 97300
rect 31076 97288 31082 97300
rect 82814 97288 82820 97300
rect 31076 97260 82820 97288
rect 31076 97248 31082 97260
rect 82814 97248 82820 97260
rect 82872 97248 82878 97300
rect 93394 97248 93400 97300
rect 93452 97288 93458 97300
rect 95050 97288 95056 97300
rect 93452 97260 95056 97288
rect 93452 97248 93458 97260
rect 95050 97248 95056 97260
rect 95108 97288 95114 97300
rect 99346 97288 99374 97328
rect 116394 97316 116400 97328
rect 116452 97316 116458 97368
rect 120074 97316 120080 97368
rect 120132 97356 120138 97368
rect 120718 97356 120724 97368
rect 120132 97328 120724 97356
rect 120132 97316 120138 97328
rect 120718 97316 120724 97328
rect 120776 97316 120782 97368
rect 295978 97356 295984 97368
rect 122852 97328 295984 97356
rect 95108 97260 99374 97288
rect 95108 97248 95114 97260
rect 104894 97248 104900 97300
rect 104952 97288 104958 97300
rect 105538 97288 105544 97300
rect 104952 97260 105544 97288
rect 104952 97248 104958 97260
rect 105538 97248 105544 97260
rect 105596 97248 105602 97300
rect 110414 97248 110420 97300
rect 110472 97288 110478 97300
rect 110472 97260 115934 97288
rect 110472 97248 110478 97260
rect 81526 97180 81532 97232
rect 81584 97220 81590 97232
rect 91002 97220 91008 97232
rect 81584 97192 91008 97220
rect 81584 97180 81590 97192
rect 91002 97180 91008 97192
rect 91060 97220 91066 97232
rect 93670 97220 93676 97232
rect 91060 97192 93676 97220
rect 91060 97180 91066 97192
rect 93670 97180 93676 97192
rect 93728 97180 93734 97232
rect 94958 97180 94964 97232
rect 95016 97220 95022 97232
rect 95016 97192 99374 97220
rect 95016 97180 95022 97192
rect 89530 97112 89536 97164
rect 89588 97152 89594 97164
rect 90450 97152 90456 97164
rect 89588 97124 90456 97152
rect 89588 97112 89594 97124
rect 90450 97112 90456 97124
rect 90508 97112 90514 97164
rect 97258 97112 97264 97164
rect 97316 97152 97322 97164
rect 97534 97152 97540 97164
rect 97316 97124 97540 97152
rect 97316 97112 97322 97124
rect 97534 97112 97540 97124
rect 97592 97112 97598 97164
rect 81802 97044 81808 97096
rect 81860 97084 81866 97096
rect 87782 97084 87788 97096
rect 81860 97056 87788 97084
rect 81860 97044 81866 97056
rect 87782 97044 87788 97056
rect 87840 97044 87846 97096
rect 91554 97044 91560 97096
rect 91612 97084 91618 97096
rect 94774 97084 94780 97096
rect 91612 97056 94780 97084
rect 91612 97044 91618 97056
rect 94774 97044 94780 97056
rect 94832 97044 94838 97096
rect 71038 96976 71044 97028
rect 71096 97016 71102 97028
rect 85482 97016 85488 97028
rect 71096 96988 85488 97016
rect 71096 96976 71102 96988
rect 85482 96976 85488 96988
rect 85540 96976 85546 97028
rect 82170 96908 82176 96960
rect 82228 96948 82234 96960
rect 82228 96920 86724 96948
rect 82228 96908 82234 96920
rect 86696 96812 86724 96920
rect 93394 96812 93400 96824
rect 86696 96784 93400 96812
rect 93394 96772 93400 96784
rect 93452 96772 93458 96824
rect 87414 96744 87420 96756
rect 86236 96716 87420 96744
rect 82630 96636 82636 96688
rect 82688 96676 82694 96688
rect 83090 96676 83096 96688
rect 82688 96648 83096 96676
rect 82688 96636 82694 96648
rect 83090 96636 83096 96648
rect 83148 96636 83154 96688
rect 85666 96568 85672 96620
rect 85724 96608 85730 96620
rect 86236 96608 86264 96716
rect 87414 96704 87420 96716
rect 87472 96704 87478 96756
rect 86402 96636 86408 96688
rect 86460 96676 86466 96688
rect 87506 96676 87512 96688
rect 86460 96648 87512 96676
rect 86460 96636 86466 96648
rect 87506 96636 87512 96648
rect 87564 96636 87570 96688
rect 92474 96636 92480 96688
rect 92532 96676 92538 96688
rect 93394 96676 93400 96688
rect 92532 96648 93400 96676
rect 92532 96636 92538 96648
rect 93394 96636 93400 96648
rect 93452 96636 93458 96688
rect 99346 96676 99374 97192
rect 110598 97112 110604 97164
rect 110656 97152 110662 97164
rect 111150 97152 111156 97164
rect 110656 97124 111156 97152
rect 110656 97112 110662 97124
rect 111150 97112 111156 97124
rect 111208 97112 111214 97164
rect 105170 96976 105176 97028
rect 105228 97016 105234 97028
rect 105446 97016 105452 97028
rect 105228 96988 105452 97016
rect 105228 96976 105234 96988
rect 105446 96976 105452 96988
rect 105504 96976 105510 97028
rect 115906 97016 115934 97260
rect 118970 97248 118976 97300
rect 119028 97288 119034 97300
rect 119614 97288 119620 97300
rect 119028 97260 119620 97288
rect 119028 97248 119034 97260
rect 119614 97248 119620 97260
rect 119672 97248 119678 97300
rect 119706 97248 119712 97300
rect 119764 97288 119770 97300
rect 122852 97288 122880 97328
rect 295978 97316 295984 97328
rect 296036 97316 296042 97368
rect 119764 97260 122880 97288
rect 119764 97248 119770 97260
rect 124490 97248 124496 97300
rect 124548 97288 124554 97300
rect 446398 97288 446404 97300
rect 124548 97260 446404 97288
rect 124548 97248 124554 97260
rect 446398 97248 446404 97260
rect 446456 97248 446462 97300
rect 118602 97180 118608 97232
rect 118660 97220 118666 97232
rect 129090 97220 129096 97232
rect 118660 97192 129096 97220
rect 118660 97180 118666 97192
rect 129090 97180 129096 97192
rect 129148 97180 129154 97232
rect 119154 97112 119160 97164
rect 119212 97152 119218 97164
rect 129274 97152 129280 97164
rect 119212 97124 129280 97152
rect 119212 97112 119218 97124
rect 129274 97112 129280 97124
rect 129332 97112 129338 97164
rect 118142 97044 118148 97096
rect 118200 97084 118206 97096
rect 119798 97084 119804 97096
rect 118200 97056 119804 97084
rect 118200 97044 118206 97056
rect 119798 97044 119804 97056
rect 119856 97044 119862 97096
rect 121086 97016 121092 97028
rect 115906 96988 121092 97016
rect 121086 96976 121092 96988
rect 121144 96976 121150 97028
rect 114922 96908 114928 96960
rect 114980 96948 114986 96960
rect 114980 96920 118280 96948
rect 114980 96908 114986 96920
rect 105170 96840 105176 96892
rect 105228 96880 105234 96892
rect 105630 96880 105636 96892
rect 105228 96852 105636 96880
rect 105228 96840 105234 96852
rect 105630 96840 105636 96852
rect 105688 96840 105694 96892
rect 118252 96880 118280 96920
rect 118786 96908 118792 96960
rect 118844 96948 118850 96960
rect 119154 96948 119160 96960
rect 118844 96920 119160 96948
rect 118844 96908 118850 96920
rect 119154 96908 119160 96920
rect 119212 96908 119218 96960
rect 120810 96908 120816 96960
rect 120868 96948 120874 96960
rect 120994 96948 121000 96960
rect 120868 96920 121000 96948
rect 120868 96908 120874 96920
rect 120994 96908 121000 96920
rect 121052 96908 121058 96960
rect 118252 96852 118556 96880
rect 118528 96824 118556 96852
rect 118878 96840 118884 96892
rect 118936 96880 118942 96892
rect 119522 96880 119528 96892
rect 118936 96852 119528 96880
rect 118936 96840 118942 96852
rect 119522 96840 119528 96852
rect 119580 96840 119586 96892
rect 111610 96772 111616 96824
rect 111668 96812 111674 96824
rect 112806 96812 112812 96824
rect 111668 96784 112812 96812
rect 111668 96772 111674 96784
rect 112806 96772 112812 96784
rect 112864 96772 112870 96824
rect 113082 96772 113088 96824
rect 113140 96812 113146 96824
rect 114922 96812 114928 96824
rect 113140 96784 114928 96812
rect 113140 96772 113146 96784
rect 114922 96772 114928 96784
rect 114980 96772 114986 96824
rect 115750 96772 115756 96824
rect 115808 96812 115814 96824
rect 117038 96812 117044 96824
rect 115808 96784 117044 96812
rect 115808 96772 115814 96784
rect 117038 96772 117044 96784
rect 117096 96772 117102 96824
rect 118510 96772 118516 96824
rect 118568 96772 118574 96824
rect 118786 96772 118792 96824
rect 118844 96812 118850 96824
rect 119430 96812 119436 96824
rect 118844 96784 119436 96812
rect 118844 96772 118850 96784
rect 119430 96772 119436 96784
rect 119488 96772 119494 96824
rect 106458 96704 106464 96756
rect 106516 96744 106522 96756
rect 107102 96744 107108 96756
rect 106516 96716 107108 96744
rect 106516 96704 106522 96716
rect 107102 96704 107108 96716
rect 107160 96704 107166 96756
rect 113818 96704 113824 96756
rect 113876 96744 113882 96756
rect 119706 96744 119712 96756
rect 113876 96716 119712 96744
rect 113876 96704 113882 96716
rect 119706 96704 119712 96716
rect 119764 96704 119770 96756
rect 120350 96704 120356 96756
rect 120408 96744 120414 96756
rect 127986 96744 127992 96756
rect 120408 96716 127992 96744
rect 120408 96704 120414 96716
rect 127986 96704 127992 96716
rect 128044 96704 128050 96756
rect 121362 96676 121368 96688
rect 99346 96648 121368 96676
rect 121362 96636 121368 96648
rect 121420 96636 121426 96688
rect 123570 96636 123576 96688
rect 123628 96676 123634 96688
rect 125134 96676 125140 96688
rect 123628 96648 125140 96676
rect 123628 96636 123634 96648
rect 125134 96636 125140 96648
rect 125192 96636 125198 96688
rect 95326 96608 95332 96620
rect 85724 96580 86264 96608
rect 89686 96580 95332 96608
rect 85724 96568 85730 96580
rect 82262 96500 82268 96552
rect 82320 96540 82326 96552
rect 89686 96540 89714 96580
rect 95326 96568 95332 96580
rect 95384 96568 95390 96620
rect 106274 96568 106280 96620
rect 106332 96608 106338 96620
rect 106734 96608 106740 96620
rect 106332 96580 106740 96608
rect 106332 96568 106338 96580
rect 106734 96568 106740 96580
rect 106792 96568 106798 96620
rect 109126 96568 109132 96620
rect 109184 96608 109190 96620
rect 110230 96608 110236 96620
rect 109184 96580 110236 96608
rect 109184 96568 109190 96580
rect 110230 96568 110236 96580
rect 110288 96568 110294 96620
rect 118878 96568 118884 96620
rect 118936 96608 118942 96620
rect 119614 96608 119620 96620
rect 118936 96580 119620 96608
rect 118936 96568 118942 96580
rect 119614 96568 119620 96580
rect 119672 96568 119678 96620
rect 128998 96608 129004 96620
rect 128326 96580 129004 96608
rect 82320 96512 89714 96540
rect 82320 96500 82326 96512
rect 103514 96500 103520 96552
rect 103572 96540 103578 96552
rect 103882 96540 103888 96552
rect 103572 96512 103888 96540
rect 103572 96500 103578 96512
rect 103882 96500 103888 96512
rect 103940 96500 103946 96552
rect 116394 96500 116400 96552
rect 116452 96540 116458 96552
rect 116854 96540 116860 96552
rect 116452 96512 116860 96540
rect 116452 96500 116458 96512
rect 116854 96500 116860 96512
rect 116912 96500 116918 96552
rect 117682 96500 117688 96552
rect 117740 96540 117746 96552
rect 127894 96540 127900 96552
rect 117740 96512 127900 96540
rect 117740 96500 117746 96512
rect 127894 96500 127900 96512
rect 127952 96500 127958 96552
rect 94866 96432 94872 96484
rect 94924 96472 94930 96484
rect 128326 96472 128354 96580
rect 128998 96568 129004 96580
rect 129056 96568 129062 96620
rect 94924 96444 128354 96472
rect 94924 96432 94930 96444
rect 81342 96364 81348 96416
rect 81400 96404 81406 96416
rect 94222 96404 94228 96416
rect 81400 96376 94228 96404
rect 81400 96364 81406 96376
rect 94222 96364 94228 96376
rect 94280 96404 94286 96416
rect 94682 96404 94688 96416
rect 94280 96376 94688 96404
rect 94280 96364 94286 96376
rect 94682 96364 94688 96376
rect 94740 96364 94746 96416
rect 101030 96364 101036 96416
rect 101088 96404 101094 96416
rect 135990 96404 135996 96416
rect 101088 96376 135996 96404
rect 101088 96364 101094 96376
rect 135990 96364 135996 96376
rect 136048 96364 136054 96416
rect 80974 96296 80980 96348
rect 81032 96336 81038 96348
rect 93762 96336 93768 96348
rect 81032 96308 93768 96336
rect 81032 96296 81038 96308
rect 93762 96296 93768 96308
rect 93820 96336 93826 96348
rect 94590 96336 94596 96348
rect 93820 96308 94596 96336
rect 93820 96296 93826 96308
rect 94590 96296 94596 96308
rect 94648 96296 94654 96348
rect 95234 96296 95240 96348
rect 95292 96336 95298 96348
rect 176654 96336 176660 96348
rect 95292 96308 176660 96336
rect 95292 96296 95298 96308
rect 176654 96296 176660 96308
rect 176712 96296 176718 96348
rect 81434 96228 81440 96280
rect 81492 96268 81498 96280
rect 96430 96268 96436 96280
rect 81492 96240 96436 96268
rect 81492 96228 81498 96240
rect 96430 96228 96436 96240
rect 96488 96228 96494 96280
rect 96614 96228 96620 96280
rect 96672 96268 96678 96280
rect 193214 96268 193220 96280
rect 96672 96240 193220 96268
rect 96672 96228 96678 96240
rect 193214 96228 193220 96240
rect 193272 96228 193278 96280
rect 82354 96160 82360 96212
rect 82412 96200 82418 96212
rect 95970 96200 95976 96212
rect 82412 96172 95976 96200
rect 82412 96160 82418 96172
rect 95970 96160 95976 96172
rect 96028 96160 96034 96212
rect 97442 96160 97448 96212
rect 97500 96200 97506 96212
rect 200114 96200 200120 96212
rect 97500 96172 200120 96200
rect 97500 96160 97506 96172
rect 200114 96160 200120 96172
rect 200172 96160 200178 96212
rect 106826 96092 106832 96144
rect 106884 96132 106890 96144
rect 106884 96104 107148 96132
rect 106884 96092 106890 96104
rect 81250 96024 81256 96076
rect 81308 96064 81314 96076
rect 93210 96064 93216 96076
rect 81308 96036 93216 96064
rect 81308 96024 81314 96036
rect 93210 96024 93216 96036
rect 93268 96024 93274 96076
rect 103514 96024 103520 96076
rect 103572 96064 103578 96076
rect 103698 96064 103704 96076
rect 103572 96036 103704 96064
rect 103572 96024 103578 96036
rect 103698 96024 103704 96036
rect 103756 96024 103762 96076
rect 106366 96024 106372 96076
rect 106424 96064 106430 96076
rect 107010 96064 107016 96076
rect 106424 96036 107016 96064
rect 106424 96024 106430 96036
rect 107010 96024 107016 96036
rect 107068 96024 107074 96076
rect 105078 95956 105084 96008
rect 105136 95996 105142 96008
rect 105722 95996 105728 96008
rect 105136 95968 105728 95996
rect 105136 95956 105142 95968
rect 105722 95956 105728 95968
rect 105780 95956 105786 96008
rect 106274 95956 106280 96008
rect 106332 95996 106338 96008
rect 106826 95996 106832 96008
rect 106332 95968 106832 95996
rect 106332 95956 106338 95968
rect 106826 95956 106832 95968
rect 106884 95956 106890 96008
rect 107010 95888 107016 95940
rect 107068 95928 107074 95940
rect 107120 95928 107148 96104
rect 107378 96092 107384 96144
rect 107436 96132 107442 96144
rect 107930 96132 107936 96144
rect 107436 96104 107936 96132
rect 107436 96092 107442 96104
rect 107930 96092 107936 96104
rect 107988 96092 107994 96144
rect 109034 96092 109040 96144
rect 109092 96132 109098 96144
rect 109494 96132 109500 96144
rect 109092 96104 109500 96132
rect 109092 96092 109098 96104
rect 109494 96092 109500 96104
rect 109552 96092 109558 96144
rect 114922 96092 114928 96144
rect 114980 96132 114986 96144
rect 115750 96132 115756 96144
rect 114980 96104 115756 96132
rect 114980 96092 114986 96104
rect 115750 96092 115756 96104
rect 115808 96092 115814 96144
rect 117498 96092 117504 96144
rect 117556 96132 117562 96144
rect 117682 96132 117688 96144
rect 117556 96104 117688 96132
rect 117556 96092 117562 96104
rect 117682 96092 117688 96104
rect 117740 96092 117746 96144
rect 122006 96092 122012 96144
rect 122064 96132 122070 96144
rect 498194 96132 498200 96144
rect 122064 96104 498200 96132
rect 122064 96092 122070 96104
rect 498194 96092 498200 96104
rect 498252 96092 498258 96144
rect 109218 96024 109224 96076
rect 109276 96064 109282 96076
rect 109862 96064 109868 96076
rect 109276 96036 109868 96064
rect 109276 96024 109282 96036
rect 109862 96024 109868 96036
rect 109920 96024 109926 96076
rect 123846 96024 123852 96076
rect 123904 96064 123910 96076
rect 514754 96064 514760 96076
rect 123904 96036 514760 96064
rect 123904 96024 123910 96036
rect 514754 96024 514760 96036
rect 514812 96024 514818 96076
rect 114922 95956 114928 96008
rect 114980 95996 114986 96008
rect 115106 95996 115112 96008
rect 114980 95968 115112 95996
rect 114980 95956 114986 95968
rect 115106 95956 115112 95968
rect 115164 95956 115170 96008
rect 125502 95956 125508 96008
rect 125560 95996 125566 96008
rect 528554 95996 528560 96008
rect 125560 95968 528560 95996
rect 125560 95956 125566 95968
rect 528554 95956 528560 95968
rect 528612 95956 528618 96008
rect 107068 95900 107148 95928
rect 107068 95888 107074 95900
rect 126514 95888 126520 95940
rect 126572 95928 126578 95940
rect 545114 95928 545120 95940
rect 126572 95900 545120 95928
rect 126572 95888 126578 95900
rect 545114 95888 545120 95900
rect 545172 95888 545178 95940
rect 81158 95820 81164 95872
rect 81216 95860 81222 95872
rect 93302 95860 93308 95872
rect 81216 95832 93308 95860
rect 81216 95820 81222 95832
rect 93302 95820 93308 95832
rect 93360 95820 93366 95872
rect 96706 95820 96712 95872
rect 96764 95860 96770 95872
rect 97166 95860 97172 95872
rect 96764 95832 97172 95860
rect 96764 95820 96770 95832
rect 97166 95820 97172 95832
rect 97224 95820 97230 95872
rect 105078 95820 105084 95872
rect 105136 95860 105142 95872
rect 105354 95860 105360 95872
rect 105136 95832 105360 95860
rect 105136 95820 105142 95832
rect 105354 95820 105360 95832
rect 105412 95820 105418 95872
rect 106274 95820 106280 95872
rect 106332 95860 106338 95872
rect 107194 95860 107200 95872
rect 106332 95832 107200 95860
rect 106332 95820 106338 95832
rect 107194 95820 107200 95832
rect 107252 95820 107258 95872
rect 81066 95752 81072 95804
rect 81124 95792 81130 95804
rect 93578 95792 93584 95804
rect 81124 95764 93584 95792
rect 81124 95752 81130 95764
rect 93578 95752 93584 95764
rect 93636 95792 93642 95804
rect 94498 95792 94504 95804
rect 93636 95764 94504 95792
rect 93636 95752 93642 95764
rect 94498 95752 94504 95764
rect 94556 95752 94562 95804
rect 103606 95752 103612 95804
rect 103664 95792 103670 95804
rect 104342 95792 104348 95804
rect 103664 95764 104348 95792
rect 103664 95752 103670 95764
rect 104342 95752 104348 95764
rect 104400 95752 104406 95804
rect 116946 95752 116952 95804
rect 117004 95792 117010 95804
rect 122466 95792 122472 95804
rect 117004 95764 122472 95792
rect 117004 95752 117010 95764
rect 122466 95752 122472 95764
rect 122524 95752 122530 95804
rect 104986 95684 104992 95736
rect 105044 95724 105050 95736
rect 105354 95724 105360 95736
rect 105044 95696 105360 95724
rect 105044 95684 105050 95696
rect 105354 95684 105360 95696
rect 105412 95684 105418 95736
rect 109402 95616 109408 95668
rect 109460 95656 109466 95668
rect 109954 95656 109960 95668
rect 109460 95628 109960 95656
rect 109460 95616 109466 95628
rect 109954 95616 109960 95628
rect 110012 95616 110018 95668
rect 102134 95548 102140 95600
rect 102192 95588 102198 95600
rect 102594 95588 102600 95600
rect 102192 95560 102600 95588
rect 102192 95548 102198 95560
rect 102594 95548 102600 95560
rect 102652 95548 102658 95600
rect 104986 95548 104992 95600
rect 105044 95588 105050 95600
rect 105170 95588 105176 95600
rect 105044 95560 105176 95588
rect 105044 95548 105050 95560
rect 105170 95548 105176 95560
rect 105228 95548 105234 95600
rect 107746 95548 107752 95600
rect 107804 95588 107810 95600
rect 108758 95588 108764 95600
rect 107804 95560 108764 95588
rect 107804 95548 107810 95560
rect 108758 95548 108764 95560
rect 108816 95548 108822 95600
rect 110506 95548 110512 95600
rect 110564 95588 110570 95600
rect 111518 95588 111524 95600
rect 110564 95560 111524 95588
rect 110564 95548 110570 95560
rect 111518 95548 111524 95560
rect 111576 95548 111582 95600
rect 102226 95412 102232 95464
rect 102284 95452 102290 95464
rect 102594 95452 102600 95464
rect 102284 95424 102600 95452
rect 102284 95412 102290 95424
rect 102594 95412 102600 95424
rect 102652 95412 102658 95464
rect 115842 95344 115848 95396
rect 115900 95384 115906 95396
rect 118142 95384 118148 95396
rect 115900 95356 118148 95384
rect 115900 95344 115906 95356
rect 118142 95344 118148 95356
rect 118200 95344 118206 95396
rect 121546 95344 121552 95396
rect 121604 95384 121610 95396
rect 121914 95384 121920 95396
rect 121604 95356 121920 95384
rect 121604 95344 121610 95356
rect 121914 95344 121920 95356
rect 121972 95344 121978 95396
rect 95326 95208 95332 95260
rect 95384 95248 95390 95260
rect 96154 95248 96160 95260
rect 95384 95220 96160 95248
rect 95384 95208 95390 95220
rect 96154 95208 96160 95220
rect 96212 95208 96218 95260
rect 114830 95140 114836 95192
rect 114888 95180 114894 95192
rect 115474 95180 115480 95192
rect 114888 95152 115480 95180
rect 114888 95140 114894 95152
rect 115474 95140 115480 95152
rect 115532 95140 115538 95192
rect 121454 95140 121460 95192
rect 121512 95180 121518 95192
rect 121822 95180 121828 95192
rect 121512 95152 121828 95180
rect 121512 95140 121518 95152
rect 121822 95140 121828 95152
rect 121880 95140 121886 95192
rect 110230 95072 110236 95124
rect 110288 95112 110294 95124
rect 115842 95112 115848 95124
rect 110288 95084 115848 95112
rect 110288 95072 110294 95084
rect 115842 95072 115848 95084
rect 115900 95072 115906 95124
rect 113450 95004 113456 95056
rect 113508 95044 113514 95056
rect 113818 95044 113824 95056
rect 113508 95016 113824 95044
rect 113508 95004 113514 95016
rect 113818 95004 113824 95016
rect 113876 95004 113882 95056
rect 116026 95004 116032 95056
rect 116084 95044 116090 95056
rect 116394 95044 116400 95056
rect 116084 95016 116400 95044
rect 116084 95004 116090 95016
rect 116394 95004 116400 95016
rect 116452 95004 116458 95056
rect 126974 95044 126980 95056
rect 118666 95016 126980 95044
rect 91278 94936 91284 94988
rect 91336 94976 91342 94988
rect 118666 94976 118694 95016
rect 126974 95004 126980 95016
rect 127032 95004 127038 95056
rect 91336 94948 118694 94976
rect 91336 94936 91342 94948
rect 121638 94936 121644 94988
rect 121696 94976 121702 94988
rect 122558 94976 122564 94988
rect 121696 94948 122564 94976
rect 121696 94936 121702 94948
rect 122558 94936 122564 94948
rect 122616 94936 122622 94988
rect 123294 94936 123300 94988
rect 123352 94976 123358 94988
rect 123478 94976 123484 94988
rect 123352 94948 123484 94976
rect 123352 94936 123358 94948
rect 123478 94936 123484 94948
rect 123536 94936 123542 94988
rect 107470 94868 107476 94920
rect 107528 94908 107534 94920
rect 162118 94908 162124 94920
rect 107528 94880 162124 94908
rect 107528 94868 107534 94880
rect 162118 94868 162124 94880
rect 162176 94868 162182 94920
rect 96614 94800 96620 94852
rect 96672 94840 96678 94852
rect 97902 94840 97908 94852
rect 96672 94812 97908 94840
rect 96672 94800 96678 94812
rect 97902 94800 97908 94812
rect 97960 94800 97966 94852
rect 101214 94800 101220 94852
rect 101272 94840 101278 94852
rect 247034 94840 247040 94852
rect 101272 94812 247040 94840
rect 101272 94800 101278 94812
rect 247034 94800 247040 94812
rect 247092 94800 247098 94852
rect 84746 94732 84752 94784
rect 84804 94772 84810 94784
rect 85114 94772 85120 94784
rect 84804 94744 85120 94772
rect 84804 94732 84810 94744
rect 85114 94732 85120 94744
rect 85172 94732 85178 94784
rect 88702 94732 88708 94784
rect 88760 94772 88766 94784
rect 89070 94772 89076 94784
rect 88760 94744 89076 94772
rect 88760 94732 88766 94744
rect 89070 94732 89076 94744
rect 89128 94732 89134 94784
rect 101858 94732 101864 94784
rect 101916 94772 101922 94784
rect 252554 94772 252560 94784
rect 101916 94744 252560 94772
rect 101916 94732 101922 94744
rect 252554 94732 252560 94744
rect 252612 94732 252618 94784
rect 81526 94664 81532 94716
rect 81584 94704 81590 94716
rect 82446 94704 82452 94716
rect 81584 94676 82452 94704
rect 81584 94664 81590 94676
rect 82446 94664 82452 94676
rect 82504 94664 82510 94716
rect 83366 94664 83372 94716
rect 83424 94704 83430 94716
rect 83642 94704 83648 94716
rect 83424 94676 83648 94704
rect 83424 94664 83430 94676
rect 83642 94664 83648 94676
rect 83700 94664 83706 94716
rect 85022 94664 85028 94716
rect 85080 94704 85086 94716
rect 85390 94704 85396 94716
rect 85080 94676 85396 94704
rect 85080 94664 85086 94676
rect 85390 94664 85396 94676
rect 85448 94664 85454 94716
rect 87138 94664 87144 94716
rect 87196 94664 87202 94716
rect 87230 94664 87236 94716
rect 87288 94704 87294 94716
rect 87506 94704 87512 94716
rect 87288 94676 87512 94704
rect 87288 94664 87294 94676
rect 87506 94664 87512 94676
rect 87564 94664 87570 94716
rect 88794 94664 88800 94716
rect 88852 94664 88858 94716
rect 95878 94664 95884 94716
rect 95936 94704 95942 94716
rect 96338 94704 96344 94716
rect 95936 94676 96344 94704
rect 95936 94664 95942 94676
rect 96338 94664 96344 94676
rect 96396 94664 96402 94716
rect 96798 94664 96804 94716
rect 96856 94664 96862 94716
rect 98086 94664 98092 94716
rect 98144 94704 98150 94716
rect 99282 94704 99288 94716
rect 98144 94676 99288 94704
rect 98144 94664 98150 94676
rect 99282 94664 99288 94676
rect 99340 94664 99346 94716
rect 103330 94664 103336 94716
rect 103388 94704 103394 94716
rect 266354 94704 266360 94716
rect 103388 94676 266360 94704
rect 103388 94664 103394 94676
rect 266354 94664 266360 94676
rect 266412 94664 266418 94716
rect 87156 94636 87184 94664
rect 87156 94608 88196 94636
rect 83090 94528 83096 94580
rect 83148 94568 83154 94580
rect 83458 94568 83464 94580
rect 83148 94540 83464 94568
rect 83148 94528 83154 94540
rect 83458 94528 83464 94540
rect 83516 94528 83522 94580
rect 85850 94528 85856 94580
rect 85908 94568 85914 94580
rect 86310 94568 86316 94580
rect 85908 94540 86316 94568
rect 85908 94528 85914 94540
rect 86310 94528 86316 94540
rect 86368 94528 86374 94580
rect 86954 94528 86960 94580
rect 87012 94568 87018 94580
rect 87598 94568 87604 94580
rect 87012 94540 87604 94568
rect 87012 94528 87018 94540
rect 87598 94528 87604 94540
rect 87656 94528 87662 94580
rect 87414 94460 87420 94512
rect 87472 94500 87478 94512
rect 88058 94500 88064 94512
rect 87472 94472 88064 94500
rect 87472 94460 87478 94472
rect 88058 94460 88064 94472
rect 88116 94460 88122 94512
rect 82906 94392 82912 94444
rect 82964 94432 82970 94444
rect 83458 94432 83464 94444
rect 82964 94404 83464 94432
rect 82964 94392 82970 94404
rect 83458 94392 83464 94404
rect 83516 94392 83522 94444
rect 83550 94392 83556 94444
rect 83608 94432 83614 94444
rect 83734 94432 83740 94444
rect 83608 94404 83740 94432
rect 83608 94392 83614 94404
rect 83734 94392 83740 94404
rect 83792 94392 83798 94444
rect 84838 94392 84844 94444
rect 84896 94432 84902 94444
rect 85298 94432 85304 94444
rect 84896 94404 85304 94432
rect 84896 94392 84902 94404
rect 85298 94392 85304 94404
rect 85356 94392 85362 94444
rect 85850 94392 85856 94444
rect 85908 94432 85914 94444
rect 86862 94432 86868 94444
rect 85908 94404 86868 94432
rect 85908 94392 85914 94404
rect 86862 94392 86868 94404
rect 86920 94392 86926 94444
rect 87138 94392 87144 94444
rect 87196 94432 87202 94444
rect 87874 94432 87880 94444
rect 87196 94404 87880 94432
rect 87196 94392 87202 94404
rect 87874 94392 87880 94404
rect 87932 94392 87938 94444
rect 84378 94324 84384 94376
rect 84436 94364 84442 94376
rect 84930 94364 84936 94376
rect 84436 94336 84936 94364
rect 84436 94324 84442 94336
rect 84930 94324 84936 94336
rect 84988 94324 84994 94376
rect 85942 94324 85948 94376
rect 86000 94364 86006 94376
rect 86770 94364 86776 94376
rect 86000 94336 86776 94364
rect 86000 94324 86006 94336
rect 86770 94324 86776 94336
rect 86828 94324 86834 94376
rect 88058 94324 88064 94376
rect 88116 94364 88122 94376
rect 88168 94364 88196 94608
rect 88334 94568 88340 94580
rect 88116 94336 88196 94364
rect 88260 94540 88340 94568
rect 88260 94364 88288 94540
rect 88334 94528 88340 94540
rect 88392 94528 88398 94580
rect 88334 94392 88340 94444
rect 88392 94432 88398 94444
rect 88812 94432 88840 94664
rect 91370 94596 91376 94648
rect 91428 94636 91434 94648
rect 91830 94636 91836 94648
rect 91428 94608 91836 94636
rect 91428 94596 91434 94608
rect 91830 94596 91836 94608
rect 91888 94596 91894 94648
rect 90082 94528 90088 94580
rect 90140 94568 90146 94580
rect 90266 94568 90272 94580
rect 90140 94540 90272 94568
rect 90140 94528 90146 94540
rect 90266 94528 90272 94540
rect 90324 94528 90330 94580
rect 91278 94528 91284 94580
rect 91336 94568 91342 94580
rect 91922 94568 91928 94580
rect 91336 94540 91928 94568
rect 91336 94528 91342 94540
rect 91922 94528 91928 94540
rect 91980 94528 91986 94580
rect 93854 94528 93860 94580
rect 93912 94568 93918 94580
rect 94038 94568 94044 94580
rect 93912 94540 94044 94568
rect 93912 94528 93918 94540
rect 94038 94528 94044 94540
rect 94096 94528 94102 94580
rect 94222 94528 94228 94580
rect 94280 94568 94286 94580
rect 94406 94568 94412 94580
rect 94280 94540 94412 94568
rect 94280 94528 94286 94540
rect 94406 94528 94412 94540
rect 94464 94528 94470 94580
rect 95510 94528 95516 94580
rect 95568 94568 95574 94580
rect 95786 94568 95792 94580
rect 95568 94540 95792 94568
rect 95568 94528 95574 94540
rect 95786 94528 95792 94540
rect 95844 94528 95850 94580
rect 95878 94528 95884 94580
rect 95936 94568 95942 94580
rect 96062 94568 96068 94580
rect 95936 94540 96068 94568
rect 95936 94528 95942 94540
rect 96062 94528 96068 94540
rect 96120 94528 96126 94580
rect 96816 94512 96844 94664
rect 97994 94596 98000 94648
rect 98052 94636 98058 94648
rect 98362 94636 98368 94648
rect 98052 94608 98368 94636
rect 98052 94596 98058 94608
rect 98362 94596 98368 94608
rect 98420 94596 98426 94648
rect 105998 94596 106004 94648
rect 106056 94636 106062 94648
rect 296714 94636 296720 94648
rect 106056 94608 296720 94636
rect 106056 94596 106062 94608
rect 296714 94596 296720 94608
rect 296772 94596 296778 94648
rect 98086 94528 98092 94580
rect 98144 94568 98150 94580
rect 98270 94568 98276 94580
rect 98144 94540 98276 94568
rect 98144 94528 98150 94540
rect 98270 94528 98276 94540
rect 98328 94528 98334 94580
rect 100018 94528 100024 94580
rect 100076 94568 100082 94580
rect 100662 94568 100668 94580
rect 100076 94540 100668 94568
rect 100076 94528 100082 94540
rect 100662 94528 100668 94540
rect 100720 94528 100726 94580
rect 100938 94528 100944 94580
rect 100996 94568 101002 94580
rect 101582 94568 101588 94580
rect 100996 94540 101588 94568
rect 100996 94528 101002 94540
rect 101582 94528 101588 94540
rect 101640 94528 101646 94580
rect 109586 94568 109592 94580
rect 108960 94540 109592 94568
rect 108960 94512 108988 94540
rect 109586 94528 109592 94540
rect 109644 94528 109650 94580
rect 111794 94528 111800 94580
rect 111852 94568 111858 94580
rect 111978 94568 111984 94580
rect 111852 94540 111984 94568
rect 111852 94528 111858 94540
rect 111978 94528 111984 94540
rect 112036 94528 112042 94580
rect 112070 94528 112076 94580
rect 112128 94568 112134 94580
rect 112128 94540 112668 94568
rect 112128 94528 112134 94540
rect 89898 94460 89904 94512
rect 89956 94500 89962 94512
rect 90634 94500 90640 94512
rect 89956 94472 90640 94500
rect 89956 94460 89962 94472
rect 90634 94460 90640 94472
rect 90692 94460 90698 94512
rect 91830 94460 91836 94512
rect 91888 94500 91894 94512
rect 92382 94500 92388 94512
rect 91888 94472 92388 94500
rect 91888 94460 91894 94472
rect 92382 94460 92388 94472
rect 92440 94460 92446 94512
rect 96798 94460 96804 94512
rect 96856 94460 96862 94512
rect 96890 94460 96896 94512
rect 96948 94500 96954 94512
rect 97350 94500 97356 94512
rect 96948 94472 97356 94500
rect 96948 94460 96954 94472
rect 97350 94460 97356 94472
rect 97408 94460 97414 94512
rect 108942 94460 108948 94512
rect 109000 94460 109006 94512
rect 88392 94404 88840 94432
rect 88392 94392 88398 94404
rect 89806 94392 89812 94444
rect 89864 94432 89870 94444
rect 90266 94432 90272 94444
rect 89864 94404 90272 94432
rect 89864 94392 89870 94404
rect 90266 94392 90272 94404
rect 90324 94392 90330 94444
rect 91094 94392 91100 94444
rect 91152 94432 91158 94444
rect 91922 94432 91928 94444
rect 91152 94404 91928 94432
rect 91152 94392 91158 94404
rect 91922 94392 91928 94404
rect 91980 94392 91986 94444
rect 93762 94392 93768 94444
rect 93820 94432 93826 94444
rect 94038 94432 94044 94444
rect 93820 94404 94044 94432
rect 93820 94392 93826 94404
rect 94038 94392 94044 94404
rect 94096 94392 94102 94444
rect 101030 94392 101036 94444
rect 101088 94432 101094 94444
rect 101214 94432 101220 94444
rect 101088 94404 101220 94432
rect 101088 94392 101094 94404
rect 101214 94392 101220 94404
rect 101272 94392 101278 94444
rect 108850 94392 108856 94444
rect 108908 94432 108914 94444
rect 109586 94432 109592 94444
rect 108908 94404 109592 94432
rect 108908 94392 108914 94404
rect 109586 94392 109592 94404
rect 109644 94392 109650 94444
rect 88518 94364 88524 94376
rect 88260 94336 88524 94364
rect 88116 94324 88122 94336
rect 88518 94324 88524 94336
rect 88576 94324 88582 94376
rect 88610 94324 88616 94376
rect 88668 94364 88674 94376
rect 89622 94364 89628 94376
rect 88668 94336 89628 94364
rect 88668 94324 88674 94336
rect 89622 94324 89628 94336
rect 89680 94324 89686 94376
rect 92566 94324 92572 94376
rect 92624 94364 92630 94376
rect 93026 94364 93032 94376
rect 92624 94336 93032 94364
rect 92624 94324 92630 94336
rect 93026 94324 93032 94336
rect 93084 94324 93090 94376
rect 95970 94324 95976 94376
rect 96028 94364 96034 94376
rect 96522 94364 96528 94376
rect 96028 94336 96528 94364
rect 96028 94324 96034 94336
rect 96522 94324 96528 94336
rect 96580 94324 96586 94376
rect 98362 94324 98368 94376
rect 98420 94364 98426 94376
rect 98730 94364 98736 94376
rect 98420 94336 98736 94364
rect 98420 94324 98426 94336
rect 98730 94324 98736 94336
rect 98788 94324 98794 94376
rect 112162 94324 112168 94376
rect 112220 94364 112226 94376
rect 112530 94364 112536 94376
rect 112220 94336 112536 94364
rect 112220 94324 112226 94336
rect 112530 94324 112536 94336
rect 112588 94324 112594 94376
rect 89806 94256 89812 94308
rect 89864 94296 89870 94308
rect 90542 94296 90548 94308
rect 89864 94268 90548 94296
rect 89864 94256 89870 94268
rect 90542 94256 90548 94268
rect 90600 94256 90606 94308
rect 97902 94256 97908 94308
rect 97960 94296 97966 94308
rect 98454 94296 98460 94308
rect 97960 94268 98460 94296
rect 97960 94256 97966 94268
rect 98454 94256 98460 94268
rect 98512 94256 98518 94308
rect 112070 94256 112076 94308
rect 112128 94296 112134 94308
rect 112438 94296 112444 94308
rect 112128 94268 112444 94296
rect 112128 94256 112134 94268
rect 112438 94256 112444 94268
rect 112496 94256 112502 94308
rect 92566 94188 92572 94240
rect 92624 94228 92630 94240
rect 93670 94228 93676 94240
rect 92624 94200 93676 94228
rect 92624 94188 92630 94200
rect 93670 94188 93676 94200
rect 93728 94188 93734 94240
rect 112530 94188 112536 94240
rect 112588 94228 112594 94240
rect 112640 94228 112668 94540
rect 116026 94528 116032 94580
rect 116084 94568 116090 94580
rect 116302 94568 116308 94580
rect 116084 94540 116308 94568
rect 116084 94528 116090 94540
rect 116302 94528 116308 94540
rect 116360 94528 116366 94580
rect 342254 94568 342260 94580
rect 118528 94540 342260 94568
rect 113542 94460 113548 94512
rect 113600 94500 113606 94512
rect 113726 94500 113732 94512
rect 113600 94472 113732 94500
rect 113600 94460 113606 94472
rect 113726 94460 113732 94472
rect 113784 94460 113790 94512
rect 115198 94460 115204 94512
rect 115256 94500 115262 94512
rect 115382 94500 115388 94512
rect 115256 94472 115388 94500
rect 115256 94460 115262 94472
rect 115382 94460 115388 94472
rect 115440 94460 115446 94512
rect 115842 94460 115848 94512
rect 115900 94500 115906 94512
rect 118528 94500 118556 94540
rect 342254 94528 342260 94540
rect 342312 94528 342318 94580
rect 398834 94500 398840 94512
rect 115900 94472 118556 94500
rect 118666 94472 398840 94500
rect 115900 94460 115906 94472
rect 113266 94392 113272 94444
rect 113324 94432 113330 94444
rect 114094 94432 114100 94444
rect 113324 94404 114100 94432
rect 113324 94392 113330 94404
rect 114094 94392 114100 94404
rect 114152 94392 114158 94444
rect 114554 94392 114560 94444
rect 114612 94432 114618 94444
rect 115106 94432 115112 94444
rect 114612 94404 115112 94432
rect 114612 94392 114618 94404
rect 115106 94392 115112 94404
rect 115164 94392 115170 94444
rect 116302 94392 116308 94444
rect 116360 94432 116366 94444
rect 116762 94432 116768 94444
rect 116360 94404 116768 94432
rect 116360 94392 116366 94404
rect 116762 94392 116768 94404
rect 116820 94392 116826 94444
rect 118326 94392 118332 94444
rect 118384 94432 118390 94444
rect 118510 94432 118516 94444
rect 118384 94404 118516 94432
rect 118384 94392 118390 94404
rect 118510 94392 118516 94404
rect 118568 94392 118574 94444
rect 113082 94324 113088 94376
rect 113140 94364 113146 94376
rect 113726 94364 113732 94376
rect 113140 94336 113732 94364
rect 113140 94324 113146 94336
rect 113726 94324 113732 94336
rect 113784 94324 113790 94376
rect 114738 94324 114744 94376
rect 114796 94364 114802 94376
rect 115566 94364 115572 94376
rect 114796 94336 115572 94364
rect 114796 94324 114802 94336
rect 115566 94324 115572 94336
rect 115624 94324 115630 94376
rect 117314 94324 117320 94376
rect 117372 94364 117378 94376
rect 117866 94364 117872 94376
rect 117372 94336 117872 94364
rect 117372 94324 117378 94336
rect 117866 94324 117872 94336
rect 117924 94324 117930 94376
rect 114462 94256 114468 94308
rect 114520 94296 114526 94308
rect 118666 94296 118694 94472
rect 398834 94460 398840 94472
rect 398892 94460 398898 94512
rect 121914 94392 121920 94444
rect 121972 94432 121978 94444
rect 122282 94432 122288 94444
rect 121972 94404 122288 94432
rect 121972 94392 121978 94404
rect 122282 94392 122288 94404
rect 122340 94392 122346 94444
rect 122926 94392 122932 94444
rect 122984 94432 122990 94444
rect 123294 94432 123300 94444
rect 122984 94404 123300 94432
rect 122984 94392 122990 94404
rect 123294 94392 123300 94404
rect 123352 94392 123358 94444
rect 124490 94392 124496 94444
rect 124548 94432 124554 94444
rect 124766 94432 124772 94444
rect 124548 94404 124772 94432
rect 124548 94392 124554 94404
rect 124766 94392 124772 94404
rect 124824 94392 124830 94444
rect 123018 94324 123024 94376
rect 123076 94364 123082 94376
rect 123386 94364 123392 94376
rect 123076 94336 123392 94364
rect 123076 94324 123082 94336
rect 123386 94324 123392 94336
rect 123444 94324 123450 94376
rect 114520 94268 118694 94296
rect 114520 94256 114526 94268
rect 121638 94256 121644 94308
rect 121696 94296 121702 94308
rect 122374 94296 122380 94308
rect 121696 94268 122380 94296
rect 121696 94256 121702 94268
rect 122374 94256 122380 94268
rect 122432 94256 122438 94308
rect 122742 94256 122748 94308
rect 122800 94296 122806 94308
rect 123294 94296 123300 94308
rect 122800 94268 123300 94296
rect 122800 94256 122806 94268
rect 123294 94256 123300 94268
rect 123352 94256 123358 94308
rect 124398 94256 124404 94308
rect 124456 94296 124462 94308
rect 124766 94296 124772 94308
rect 124456 94268 124772 94296
rect 124456 94256 124462 94268
rect 124766 94256 124772 94268
rect 124824 94256 124830 94308
rect 112588 94200 112668 94228
rect 112588 94188 112594 94200
rect 123018 94188 123024 94240
rect 123076 94228 123082 94240
rect 123754 94228 123760 94240
rect 123076 94200 123760 94228
rect 123076 94188 123082 94200
rect 123754 94188 123760 94200
rect 123812 94188 123818 94240
rect 107838 94120 107844 94172
rect 107896 94160 107902 94172
rect 108482 94160 108488 94172
rect 107896 94132 108488 94160
rect 107896 94120 107902 94132
rect 108482 94120 108488 94132
rect 108540 94120 108546 94172
rect 111702 94120 111708 94172
rect 111760 94160 111766 94172
rect 112438 94160 112444 94172
rect 111760 94132 112444 94160
rect 111760 94120 111766 94132
rect 112438 94120 112444 94132
rect 112496 94120 112502 94172
rect 120166 94120 120172 94172
rect 120224 94160 120230 94172
rect 121270 94160 121276 94172
rect 120224 94132 121276 94160
rect 120224 94120 120230 94132
rect 121270 94120 121276 94132
rect 121328 94120 121334 94172
rect 124398 94120 124404 94172
rect 124456 94160 124462 94172
rect 125042 94160 125048 94172
rect 124456 94132 125048 94160
rect 124456 94120 124462 94132
rect 125042 94120 125048 94132
rect 125100 94120 125106 94172
rect 107838 93984 107844 94036
rect 107896 94024 107902 94036
rect 108206 94024 108212 94036
rect 107896 93996 108212 94024
rect 107896 93984 107902 93996
rect 108206 93984 108212 93996
rect 108264 93984 108270 94036
rect 105170 93916 105176 93968
rect 105228 93956 105234 93968
rect 105906 93956 105912 93968
rect 105228 93928 105912 93956
rect 105228 93916 105234 93928
rect 105906 93916 105912 93928
rect 105964 93916 105970 93968
rect 119522 93780 119528 93832
rect 119580 93820 119586 93832
rect 128078 93820 128084 93832
rect 119580 93792 128084 93820
rect 119580 93780 119586 93792
rect 128078 93780 128084 93792
rect 128136 93780 128142 93832
rect 110322 93712 110328 93764
rect 110380 93752 110386 93764
rect 111518 93752 111524 93764
rect 110380 93724 111524 93752
rect 110380 93712 110386 93724
rect 111518 93712 111524 93724
rect 111576 93712 111582 93764
rect 108022 93440 108028 93492
rect 108080 93480 108086 93492
rect 329834 93480 329840 93492
rect 108080 93452 329840 93480
rect 108080 93440 108086 93452
rect 329834 93440 329840 93452
rect 329892 93440 329898 93492
rect 111334 93372 111340 93424
rect 111392 93412 111398 93424
rect 346394 93412 346400 93424
rect 111392 93384 346400 93412
rect 111392 93372 111398 93384
rect 346394 93372 346400 93384
rect 346452 93372 346458 93424
rect 109770 93304 109776 93356
rect 109828 93344 109834 93356
rect 349154 93344 349160 93356
rect 109828 93316 349160 93344
rect 109828 93304 109834 93316
rect 349154 93304 349160 93316
rect 349212 93304 349218 93356
rect 112806 93236 112812 93288
rect 112864 93276 112870 93288
rect 373994 93276 374000 93288
rect 112864 93248 374000 93276
rect 112864 93236 112870 93248
rect 373994 93236 374000 93248
rect 374052 93236 374058 93288
rect 114370 93168 114376 93220
rect 114428 93208 114434 93220
rect 391934 93208 391940 93220
rect 114428 93180 391940 93208
rect 114428 93168 114434 93180
rect 391934 93168 391940 93180
rect 391992 93168 391998 93220
rect 115750 93100 115756 93152
rect 115808 93140 115814 93152
rect 401594 93140 401600 93152
rect 115808 93112 401600 93140
rect 115808 93100 115814 93112
rect 401594 93100 401600 93112
rect 401652 93100 401658 93152
rect 103422 92760 103428 92812
rect 103480 92800 103486 92812
rect 104250 92800 104256 92812
rect 103480 92772 104256 92800
rect 103480 92760 103486 92772
rect 104250 92760 104256 92772
rect 104308 92760 104314 92812
rect 101030 92488 101036 92540
rect 101088 92528 101094 92540
rect 101674 92528 101680 92540
rect 101088 92500 101680 92528
rect 101088 92488 101094 92500
rect 101674 92488 101680 92500
rect 101732 92488 101738 92540
rect 97258 92420 97264 92472
rect 97316 92460 97322 92472
rect 128814 92460 128820 92472
rect 97316 92432 128820 92460
rect 97316 92420 97322 92432
rect 128814 92420 128820 92432
rect 128872 92420 128878 92472
rect 93394 92352 93400 92404
rect 93452 92392 93458 92404
rect 142154 92392 142160 92404
rect 93452 92364 142160 92392
rect 93452 92352 93458 92364
rect 142154 92352 142160 92364
rect 142212 92352 142218 92404
rect 121362 92284 121368 92336
rect 121420 92324 121426 92336
rect 171134 92324 171140 92336
rect 121420 92296 171140 92324
rect 121420 92284 121426 92296
rect 171134 92284 171140 92296
rect 171192 92284 171198 92336
rect 116854 92216 116860 92268
rect 116912 92256 116918 92268
rect 175274 92256 175280 92268
rect 116912 92228 175280 92256
rect 116912 92216 116918 92228
rect 175274 92216 175280 92228
rect 175332 92216 175338 92268
rect 97166 92148 97172 92200
rect 97224 92188 97230 92200
rect 125042 92188 125048 92200
rect 97224 92160 125048 92188
rect 97224 92148 97230 92160
rect 125042 92148 125048 92160
rect 125100 92148 125106 92200
rect 128814 92148 128820 92200
rect 128872 92188 128878 92200
rect 194594 92188 194600 92200
rect 128872 92160 194600 92188
rect 128872 92148 128878 92160
rect 194594 92148 194600 92160
rect 194652 92148 194658 92200
rect 99466 92080 99472 92132
rect 99524 92120 99530 92132
rect 128906 92120 128912 92132
rect 99524 92092 128912 92120
rect 99524 92080 99530 92092
rect 128906 92080 128912 92092
rect 128964 92120 128970 92132
rect 224954 92120 224960 92132
rect 128964 92092 224960 92120
rect 128964 92080 128970 92092
rect 224954 92080 224960 92092
rect 225012 92080 225018 92132
rect 121086 92012 121092 92064
rect 121144 92052 121150 92064
rect 357434 92052 357440 92064
rect 121144 92024 357440 92052
rect 121144 92012 121150 92024
rect 357434 92012 357440 92024
rect 357492 92012 357498 92064
rect 114278 91944 114284 91996
rect 114336 91984 114342 91996
rect 362954 91984 362960 91996
rect 114336 91956 362960 91984
rect 114336 91944 114342 91956
rect 362954 91944 362960 91956
rect 363012 91944 363018 91996
rect 118602 91876 118608 91928
rect 118660 91916 118666 91928
rect 445754 91916 445760 91928
rect 118660 91888 445760 91916
rect 118660 91876 118666 91888
rect 445754 91876 445760 91888
rect 445812 91876 445818 91928
rect 119338 91808 119344 91860
rect 119396 91848 119402 91860
rect 456794 91848 456800 91860
rect 119396 91820 456800 91848
rect 119396 91808 119402 91820
rect 456794 91808 456800 91820
rect 456852 91808 456858 91860
rect 90358 91740 90364 91792
rect 90416 91780 90422 91792
rect 120258 91780 120264 91792
rect 90416 91752 120264 91780
rect 90416 91740 90422 91752
rect 120258 91740 120264 91752
rect 120316 91740 120322 91792
rect 125134 91740 125140 91792
rect 125192 91780 125198 91792
rect 506474 91780 506480 91792
rect 125192 91752 506480 91780
rect 125192 91740 125198 91752
rect 506474 91740 506480 91752
rect 506532 91740 506538 91792
rect 125042 91060 125048 91112
rect 125100 91100 125106 91112
rect 191834 91100 191840 91112
rect 125100 91072 191840 91100
rect 125100 91060 125106 91072
rect 191834 91060 191840 91072
rect 191892 91060 191898 91112
rect 98822 90992 98828 91044
rect 98880 91032 98886 91044
rect 128722 91032 128728 91044
rect 98880 91004 128728 91032
rect 98880 90992 98886 91004
rect 128722 90992 128728 91004
rect 128780 90992 128786 91044
rect 94590 90652 94596 90704
rect 94648 90692 94654 90704
rect 158714 90692 158720 90704
rect 94648 90664 158720 90692
rect 94648 90652 94654 90664
rect 158714 90652 158720 90664
rect 158772 90652 158778 90704
rect 128722 90584 128728 90636
rect 128780 90624 128786 90636
rect 211154 90624 211160 90636
rect 128780 90596 211160 90624
rect 128780 90584 128786 90596
rect 211154 90584 211160 90596
rect 211212 90584 211218 90636
rect 119706 90516 119712 90568
rect 119764 90556 119770 90568
rect 291194 90556 291200 90568
rect 119764 90528 291200 90556
rect 119764 90516 119770 90528
rect 291194 90516 291200 90528
rect 291252 90516 291258 90568
rect 113910 90448 113916 90500
rect 113968 90488 113974 90500
rect 307754 90488 307760 90500
rect 113968 90460 307760 90488
rect 113968 90448 113974 90460
rect 307754 90448 307760 90460
rect 307812 90448 307818 90500
rect 107102 90380 107108 90432
rect 107160 90420 107166 90432
rect 310514 90420 310520 90432
rect 107160 90392 310520 90420
rect 107160 90380 107166 90392
rect 310514 90380 310520 90392
rect 310572 90380 310578 90432
rect 91462 90312 91468 90364
rect 91520 90352 91526 90364
rect 119338 90352 119344 90364
rect 91520 90324 119344 90352
rect 91520 90312 91526 90324
rect 119338 90312 119344 90324
rect 119396 90312 119402 90364
rect 120902 90312 120908 90364
rect 120960 90352 120966 90364
rect 473446 90352 473452 90364
rect 120960 90324 473452 90352
rect 120960 90312 120966 90324
rect 473446 90312 473452 90324
rect 473504 90312 473510 90364
rect 107930 90244 107936 90296
rect 107988 90284 107994 90296
rect 108298 90284 108304 90296
rect 107988 90256 108304 90284
rect 107988 90244 107994 90256
rect 108298 90244 108304 90256
rect 108356 90244 108362 90296
rect 108022 90176 108028 90228
rect 108080 90216 108086 90228
rect 108574 90216 108580 90228
rect 108080 90188 108580 90216
rect 108080 90176 108086 90188
rect 108574 90176 108580 90188
rect 108632 90176 108638 90228
rect 102410 90108 102416 90160
rect 102468 90148 102474 90160
rect 102962 90148 102968 90160
rect 102468 90120 102968 90148
rect 102468 90108 102474 90120
rect 102962 90108 102968 90120
rect 103020 90108 103026 90160
rect 108298 90108 108304 90160
rect 108356 90148 108362 90160
rect 108482 90148 108488 90160
rect 108356 90120 108488 90148
rect 108356 90108 108362 90120
rect 108482 90108 108488 90120
rect 108540 90108 108546 90160
rect 114554 89972 114560 90024
rect 114612 90012 114618 90024
rect 115658 90012 115664 90024
rect 114612 89984 115664 90012
rect 114612 89972 114618 89984
rect 115658 89972 115664 89984
rect 115716 89972 115722 90024
rect 98546 89632 98552 89684
rect 98604 89672 98610 89684
rect 128354 89672 128360 89684
rect 98604 89644 128360 89672
rect 98604 89632 98610 89644
rect 128354 89632 128360 89644
rect 128412 89632 128418 89684
rect 92566 89564 92572 89616
rect 92624 89604 92630 89616
rect 144914 89604 144920 89616
rect 92624 89576 144920 89604
rect 92624 89564 92630 89576
rect 144914 89564 144920 89576
rect 144972 89564 144978 89616
rect 96154 89496 96160 89548
rect 96212 89536 96218 89548
rect 178034 89536 178040 89548
rect 96212 89508 178040 89536
rect 96212 89496 96218 89508
rect 178034 89496 178040 89508
rect 178092 89496 178098 89548
rect 95878 89428 95884 89480
rect 95936 89468 95942 89480
rect 180794 89468 180800 89480
rect 95936 89440 180800 89468
rect 95936 89428 95942 89440
rect 180794 89428 180800 89440
rect 180852 89428 180858 89480
rect 128354 89360 128360 89412
rect 128412 89400 128418 89412
rect 128630 89400 128636 89412
rect 128412 89372 128636 89400
rect 128412 89360 128418 89372
rect 128630 89360 128636 89372
rect 128688 89400 128694 89412
rect 218054 89400 218060 89412
rect 128688 89372 218060 89400
rect 128688 89360 128694 89372
rect 218054 89360 218060 89372
rect 218112 89360 218118 89412
rect 119798 89292 119804 89344
rect 119856 89332 119862 89344
rect 129826 89332 129832 89344
rect 119856 89304 129832 89332
rect 119856 89292 119862 89304
rect 129826 89292 129832 89304
rect 129884 89332 129890 89344
rect 241514 89332 241520 89344
rect 129884 89304 241520 89332
rect 129884 89292 129890 89304
rect 241514 89292 241520 89304
rect 241572 89292 241578 89344
rect 103238 89224 103244 89276
rect 103296 89264 103302 89276
rect 258074 89264 258080 89276
rect 103296 89236 258080 89264
rect 103296 89224 103302 89236
rect 258074 89224 258080 89236
rect 258132 89224 258138 89276
rect 104526 89156 104532 89208
rect 104584 89196 104590 89208
rect 287054 89196 287060 89208
rect 104584 89168 287060 89196
rect 104584 89156 104590 89168
rect 287054 89156 287060 89168
rect 287112 89156 287118 89208
rect 105722 89088 105728 89140
rect 105780 89128 105786 89140
rect 293954 89128 293960 89140
rect 105780 89100 293960 89128
rect 105780 89088 105786 89100
rect 293954 89088 293960 89100
rect 294012 89088 294018 89140
rect 115382 89020 115388 89072
rect 115440 89060 115446 89072
rect 409874 89060 409880 89072
rect 115440 89032 409880 89060
rect 115440 89020 115446 89032
rect 409874 89020 409880 89032
rect 409932 89020 409938 89072
rect 116670 88952 116676 89004
rect 116728 88992 116734 89004
rect 429194 88992 429200 89004
rect 116728 88964 429200 88992
rect 116728 88952 116734 88964
rect 429194 88952 429200 88964
rect 429252 88952 429258 89004
rect 127250 88884 127256 88936
rect 127308 88924 127314 88936
rect 127526 88924 127532 88936
rect 127308 88896 127532 88924
rect 127308 88884 127314 88896
rect 127526 88884 127532 88896
rect 127584 88884 127590 88936
rect 98454 88272 98460 88324
rect 98512 88312 98518 88324
rect 128446 88312 128452 88324
rect 98512 88284 128452 88312
rect 98512 88272 98518 88284
rect 128446 88272 128452 88284
rect 128504 88312 128510 88324
rect 208394 88312 208400 88324
rect 128504 88284 208400 88312
rect 128504 88272 128510 88284
rect 208394 88272 208400 88284
rect 208452 88272 208458 88324
rect 99926 88204 99932 88256
rect 99984 88244 99990 88256
rect 128538 88244 128544 88256
rect 99984 88216 128544 88244
rect 99984 88204 99990 88216
rect 128538 88204 128544 88216
rect 128596 88244 128602 88256
rect 227714 88244 227720 88256
rect 128596 88216 227720 88244
rect 128596 88204 128602 88216
rect 227714 88204 227720 88216
rect 227772 88204 227778 88256
rect 101490 88136 101496 88188
rect 101548 88176 101554 88188
rect 251174 88176 251180 88188
rect 101548 88148 251180 88176
rect 101548 88136 101554 88148
rect 251174 88136 251180 88148
rect 251232 88136 251238 88188
rect 111150 88068 111156 88120
rect 111208 88108 111214 88120
rect 360194 88108 360200 88120
rect 111208 88080 360200 88108
rect 111208 88068 111214 88080
rect 360194 88068 360200 88080
rect 360252 88068 360258 88120
rect 200758 88000 200764 88052
rect 200816 88040 200822 88052
rect 469214 88040 469220 88052
rect 200816 88012 469220 88040
rect 200816 88000 200822 88012
rect 469214 88000 469220 88012
rect 469272 88000 469278 88052
rect 115290 87932 115296 87984
rect 115348 87972 115354 87984
rect 407114 87972 407120 87984
rect 115348 87944 407120 87972
rect 115348 87932 115354 87944
rect 407114 87932 407120 87944
rect 407172 87932 407178 87984
rect 118418 87864 118424 87916
rect 118476 87904 118482 87916
rect 429286 87904 429292 87916
rect 118476 87876 429292 87904
rect 118476 87864 118482 87876
rect 429286 87864 429292 87876
rect 429344 87864 429350 87916
rect 123570 87796 123576 87848
rect 123628 87836 123634 87848
rect 511994 87836 512000 87848
rect 123628 87808 512000 87836
rect 123628 87796 123634 87808
rect 511994 87796 512000 87808
rect 512052 87796 512058 87848
rect 77294 87728 77300 87780
rect 77352 87768 77358 87780
rect 88058 87768 88064 87780
rect 77352 87740 88064 87768
rect 77352 87728 77358 87740
rect 88058 87728 88064 87740
rect 88116 87728 88122 87780
rect 123662 87728 123668 87780
rect 123720 87768 123726 87780
rect 516134 87768 516140 87780
rect 123720 87740 516140 87768
rect 123720 87728 123726 87740
rect 516134 87728 516140 87740
rect 516192 87728 516198 87780
rect 56594 87660 56600 87712
rect 56652 87700 56658 87712
rect 85482 87700 85488 87712
rect 56652 87672 85488 87700
rect 56652 87660 56658 87672
rect 85482 87660 85488 87672
rect 85540 87660 85546 87712
rect 126422 87660 126428 87712
rect 126480 87700 126486 87712
rect 545206 87700 545212 87712
rect 126480 87672 545212 87700
rect 126480 87660 126486 87672
rect 545206 87660 545212 87672
rect 545264 87660 545270 87712
rect 40034 87592 40040 87644
rect 40092 87632 40098 87644
rect 84010 87632 84016 87644
rect 40092 87604 84016 87632
rect 40092 87592 40098 87604
rect 84010 87592 84016 87604
rect 84068 87592 84074 87644
rect 91370 87592 91376 87644
rect 91428 87632 91434 87644
rect 115382 87632 115388 87644
rect 91428 87604 115388 87632
rect 91428 87592 91434 87604
rect 115382 87592 115388 87604
rect 115440 87592 115446 87644
rect 126330 87592 126336 87644
rect 126388 87632 126394 87644
rect 549254 87632 549260 87644
rect 126388 87604 549260 87632
rect 126388 87592 126394 87604
rect 549254 87592 549260 87604
rect 549312 87592 549318 87644
rect 101398 86572 101404 86624
rect 101456 86612 101462 86624
rect 244274 86612 244280 86624
rect 101456 86584 244280 86612
rect 101456 86572 101462 86584
rect 244274 86572 244280 86584
rect 244332 86572 244338 86624
rect 101306 86504 101312 86556
rect 101364 86544 101370 86556
rect 247126 86544 247132 86556
rect 101364 86516 247132 86544
rect 101364 86504 101370 86516
rect 247126 86504 247132 86516
rect 247184 86504 247190 86556
rect 104250 86436 104256 86488
rect 104308 86476 104314 86488
rect 274634 86476 274640 86488
rect 104308 86448 274640 86476
rect 104308 86436 104314 86448
rect 274634 86436 274640 86448
rect 274692 86436 274698 86488
rect 104342 86368 104348 86420
rect 104400 86408 104406 86420
rect 282914 86408 282920 86420
rect 104400 86380 282920 86408
rect 104400 86368 104406 86380
rect 282914 86368 282920 86380
rect 282972 86368 282978 86420
rect 116578 86300 116584 86352
rect 116636 86340 116642 86352
rect 433334 86340 433340 86352
rect 116636 86312 433340 86340
rect 116636 86300 116642 86312
rect 433334 86300 433340 86312
rect 433392 86300 433398 86352
rect 53834 86232 53840 86284
rect 53892 86272 53898 86284
rect 85206 86272 85212 86284
rect 53892 86244 85212 86272
rect 53892 86232 53898 86244
rect 85206 86232 85212 86244
rect 85264 86232 85270 86284
rect 117774 86232 117780 86284
rect 117832 86272 117838 86284
rect 445846 86272 445852 86284
rect 117832 86244 445852 86272
rect 117832 86232 117838 86244
rect 445846 86232 445852 86244
rect 445904 86232 445910 86284
rect 97074 85484 97080 85536
rect 97132 85524 97138 85536
rect 128354 85524 128360 85536
rect 97132 85496 128360 85524
rect 97132 85484 97138 85496
rect 128354 85484 128360 85496
rect 128412 85524 128418 85536
rect 128412 85496 132494 85524
rect 128412 85484 128418 85496
rect 132466 85252 132494 85496
rect 197354 85252 197360 85264
rect 132466 85224 197360 85252
rect 197354 85212 197360 85224
rect 197412 85212 197418 85264
rect 94314 85144 94320 85196
rect 94372 85184 94378 85196
rect 164234 85184 164240 85196
rect 94372 85156 164240 85184
rect 94372 85144 94378 85156
rect 164234 85144 164240 85156
rect 164292 85144 164298 85196
rect 108758 85076 108764 85128
rect 108816 85116 108822 85128
rect 324314 85116 324320 85128
rect 108816 85088 324320 85116
rect 108816 85076 108822 85088
rect 324314 85076 324320 85088
rect 324372 85076 324378 85128
rect 112530 85008 112536 85060
rect 112588 85048 112594 85060
rect 376754 85048 376760 85060
rect 112588 85020 376760 85048
rect 112588 85008 112594 85020
rect 376754 85008 376760 85020
rect 376812 85008 376818 85060
rect 112622 84940 112628 84992
rect 112680 84980 112686 84992
rect 379514 84980 379520 84992
rect 112680 84952 379520 84980
rect 112680 84940 112686 84952
rect 379514 84940 379520 84952
rect 379572 84940 379578 84992
rect 31754 84872 31760 84924
rect 31812 84912 31818 84924
rect 83918 84912 83924 84924
rect 31812 84884 83924 84912
rect 31812 84872 31818 84884
rect 83918 84872 83924 84884
rect 83976 84872 83982 84924
rect 116486 84872 116492 84924
rect 116544 84912 116550 84924
rect 426434 84912 426440 84924
rect 116544 84884 426440 84912
rect 116544 84872 116550 84884
rect 426434 84872 426440 84884
rect 426492 84872 426498 84924
rect 117682 84804 117688 84856
rect 117740 84844 117746 84856
rect 440234 84844 440240 84856
rect 117740 84816 440240 84844
rect 117740 84804 117746 84816
rect 440234 84804 440240 84816
rect 440292 84804 440298 84856
rect 83550 84192 83556 84244
rect 83608 84232 83614 84244
rect 86402 84232 86408 84244
rect 83608 84204 86408 84232
rect 83608 84192 83614 84204
rect 86402 84192 86408 84204
rect 86460 84192 86466 84244
rect 75914 83444 75920 83496
rect 75972 83484 75978 83496
rect 85574 83484 85580 83496
rect 75972 83456 85580 83484
rect 75972 83444 75978 83456
rect 85574 83444 85580 83456
rect 85632 83444 85638 83496
rect 109678 83444 109684 83496
rect 109736 83484 109742 83496
rect 345014 83484 345020 83496
rect 109736 83456 345020 83484
rect 109736 83444 109742 83456
rect 345014 83444 345020 83456
rect 345072 83444 345078 83496
rect 100294 82288 100300 82340
rect 100352 82328 100358 82340
rect 100570 82328 100576 82340
rect 100352 82300 100576 82328
rect 100352 82288 100358 82300
rect 100570 82288 100576 82300
rect 100628 82288 100634 82340
rect 107010 82220 107016 82272
rect 107068 82260 107074 82272
rect 313274 82260 313280 82272
rect 107068 82232 313280 82260
rect 107068 82220 107074 82232
rect 313274 82220 313280 82232
rect 313332 82220 313338 82272
rect 113818 82152 113824 82204
rect 113876 82192 113882 82204
rect 390554 82192 390560 82204
rect 113876 82164 390560 82192
rect 113876 82152 113882 82164
rect 390554 82152 390560 82164
rect 390612 82152 390618 82204
rect 123478 82084 123484 82136
rect 123536 82124 123542 82136
rect 512086 82124 512092 82136
rect 123536 82096 512092 82124
rect 123536 82084 123542 82096
rect 512086 82084 512092 82096
rect 512144 82084 512150 82136
rect 122466 80724 122472 80776
rect 122524 80764 122530 80776
rect 434714 80764 434720 80776
rect 122524 80736 434720 80764
rect 122524 80724 122530 80736
rect 434714 80724 434720 80736
rect 434772 80724 434778 80776
rect 123386 80656 123392 80708
rect 123444 80696 123450 80708
rect 507854 80696 507860 80708
rect 123444 80668 507860 80696
rect 123444 80656 123450 80668
rect 507854 80656 507860 80668
rect 507912 80656 507918 80708
rect 136082 71680 136088 71732
rect 136140 71720 136146 71732
rect 579614 71720 579620 71732
rect 136140 71692 579620 71720
rect 136140 71680 136146 71692
rect 579614 71680 579620 71692
rect 579672 71680 579678 71732
rect 129274 54476 129280 54528
rect 129332 54516 129338 54528
rect 462314 54516 462320 54528
rect 129332 54488 462320 54516
rect 129332 54476 129338 54488
rect 462314 54476 462320 54488
rect 462372 54476 462378 54528
rect 129182 53116 129188 53168
rect 129240 53156 129246 53168
rect 448514 53156 448520 53168
rect 129240 53128 448520 53156
rect 129240 53116 129246 53128
rect 448514 53116 448520 53128
rect 448572 53116 448578 53168
rect 129090 53048 129096 53100
rect 129148 53088 129154 53100
rect 455414 53088 455420 53100
rect 129148 53060 455420 53088
rect 129148 53048 129154 53060
rect 455414 53048 455420 53060
rect 455472 53048 455478 53100
rect 89162 46248 89168 46300
rect 89220 46288 89226 46300
rect 100018 46288 100024 46300
rect 89220 46260 100024 46288
rect 89220 46248 89226 46260
rect 100018 46248 100024 46260
rect 100076 46248 100082 46300
rect 99834 46180 99840 46232
rect 99892 46220 99898 46232
rect 225046 46220 225052 46232
rect 99892 46192 225052 46220
rect 99892 46180 99898 46192
rect 225046 46180 225052 46192
rect 225104 46180 225110 46232
rect 70394 44956 70400 45008
rect 70452 44996 70458 45008
rect 82630 44996 82636 45008
rect 70452 44968 82636 44996
rect 70452 44956 70458 44968
rect 82630 44956 82636 44968
rect 82688 44956 82694 45008
rect 46934 44888 46940 44940
rect 46992 44928 46998 44940
rect 84746 44928 84752 44940
rect 46992 44900 84752 44928
rect 46992 44888 46998 44900
rect 84746 44888 84752 44900
rect 84804 44888 84810 44940
rect 30374 44820 30380 44872
rect 30432 44860 30438 44872
rect 82538 44860 82544 44872
rect 30432 44832 82544 44860
rect 30432 44820 30438 44832
rect 82538 44820 82544 44832
rect 82596 44820 82602 44872
rect 94774 42100 94780 42152
rect 94832 42140 94838 42152
rect 131206 42140 131212 42152
rect 94832 42112 131212 42140
rect 94832 42100 94838 42112
rect 131206 42100 131212 42112
rect 131264 42100 131270 42152
rect 91278 42032 91284 42084
rect 91336 42072 91342 42084
rect 136726 42072 136732 42084
rect 91336 42044 136732 42072
rect 91336 42032 91342 42044
rect 136726 42032 136732 42044
rect 136784 42032 136790 42084
rect 94222 41148 94228 41200
rect 94280 41188 94286 41200
rect 165614 41188 165620 41200
rect 94280 41160 165620 41188
rect 94280 41148 94286 41160
rect 165614 41148 165620 41160
rect 165672 41148 165678 41200
rect 101214 41080 101220 41132
rect 101272 41120 101278 41132
rect 242894 41120 242900 41132
rect 101272 41092 242900 41120
rect 101272 41080 101278 41092
rect 242894 41080 242900 41092
rect 242952 41080 242958 41132
rect 105630 41012 105636 41064
rect 105688 41052 105694 41064
rect 302234 41052 302240 41064
rect 105688 41024 302240 41052
rect 105688 41012 105694 41024
rect 302234 41012 302240 41024
rect 302292 41012 302298 41064
rect 105538 40944 105544 40996
rect 105596 40984 105602 40996
rect 302326 40984 302332 40996
rect 105596 40956 302332 40984
rect 105596 40944 105602 40956
rect 302326 40944 302332 40956
rect 302384 40944 302390 40996
rect 116394 40876 116400 40928
rect 116452 40916 116458 40928
rect 423674 40916 423680 40928
rect 116452 40888 423680 40916
rect 116452 40876 116458 40888
rect 423674 40876 423680 40888
rect 423732 40876 423738 40928
rect 119154 40808 119160 40860
rect 119212 40848 119218 40860
rect 456886 40848 456892 40860
rect 119212 40820 456892 40848
rect 119212 40808 119218 40820
rect 456886 40808 456892 40820
rect 456944 40808 456950 40860
rect 119062 40740 119068 40792
rect 119120 40780 119126 40792
rect 460934 40780 460940 40792
rect 119120 40752 460940 40780
rect 119120 40740 119126 40752
rect 460934 40740 460940 40752
rect 460992 40740 460998 40792
rect 119246 40672 119252 40724
rect 119304 40712 119310 40724
rect 465074 40712 465080 40724
rect 119304 40684 465080 40712
rect 119304 40672 119310 40684
rect 465074 40672 465080 40684
rect 465132 40672 465138 40724
rect 100478 39720 100484 39772
rect 100536 39760 100542 39772
rect 237374 39760 237380 39772
rect 100536 39732 237380 39760
rect 100536 39720 100542 39732
rect 237374 39720 237380 39732
rect 237432 39720 237438 39772
rect 109586 39652 109592 39704
rect 109644 39692 109650 39704
rect 340874 39692 340880 39704
rect 109644 39664 340880 39692
rect 109644 39652 109650 39664
rect 340874 39652 340880 39664
rect 340932 39652 340938 39704
rect 112438 39584 112444 39636
rect 112496 39624 112502 39636
rect 374086 39624 374092 39636
rect 112496 39596 374092 39624
rect 112496 39584 112502 39596
rect 374086 39584 374092 39596
rect 374144 39584 374150 39636
rect 117590 39516 117596 39568
rect 117648 39556 117654 39568
rect 442994 39556 443000 39568
rect 117648 39528 443000 39556
rect 117648 39516 117654 39528
rect 442994 39516 443000 39528
rect 443052 39516 443058 39568
rect 120810 39448 120816 39500
rect 120868 39488 120874 39500
rect 483014 39488 483020 39500
rect 120868 39460 483020 39488
rect 120868 39448 120874 39460
rect 483014 39448 483020 39460
rect 483072 39448 483078 39500
rect 124950 39380 124956 39432
rect 125008 39420 125014 39432
rect 532694 39420 532700 39432
rect 125008 39392 532700 39420
rect 125008 39380 125014 39392
rect 532694 39380 532700 39392
rect 532752 39380 532758 39432
rect 126238 39312 126244 39364
rect 126296 39352 126302 39364
rect 542354 39352 542360 39364
rect 126296 39324 542360 39352
rect 126296 39312 126302 39324
rect 542354 39312 542360 39324
rect 542412 39312 542418 39364
rect 99650 38224 99656 38276
rect 99708 38264 99714 38276
rect 230474 38264 230480 38276
rect 99708 38236 230480 38264
rect 99708 38224 99714 38236
rect 230474 38224 230480 38236
rect 230532 38224 230538 38276
rect 99742 38156 99748 38208
rect 99800 38196 99806 38208
rect 233234 38196 233240 38208
rect 99800 38168 233240 38196
rect 99800 38156 99806 38168
rect 233234 38156 233240 38168
rect 233292 38156 233298 38208
rect 118326 38088 118332 38140
rect 118384 38128 118390 38140
rect 415394 38128 415400 38140
rect 118384 38100 415400 38128
rect 118384 38088 118390 38100
rect 415394 38088 415400 38100
rect 415452 38088 415458 38140
rect 116946 38020 116952 38072
rect 117004 38060 117010 38072
rect 422294 38060 422300 38072
rect 117004 38032 422300 38060
rect 117004 38020 117010 38032
rect 422294 38020 422300 38032
rect 422352 38020 422358 38072
rect 116210 37952 116216 38004
rect 116268 37992 116274 38004
rect 425054 37992 425060 38004
rect 116268 37964 425060 37992
rect 116268 37952 116274 37964
rect 425054 37952 425060 37964
rect 425112 37952 425118 38004
rect 116302 37884 116308 37936
rect 116360 37924 116366 37936
rect 431954 37924 431960 37936
rect 116360 37896 431960 37924
rect 116360 37884 116366 37896
rect 431954 37884 431960 37896
rect 432012 37884 432018 37936
rect 95694 36660 95700 36712
rect 95752 36700 95758 36712
rect 180886 36700 180892 36712
rect 95752 36672 180892 36700
rect 95752 36660 95758 36672
rect 180886 36660 180892 36672
rect 180944 36660 180950 36712
rect 96982 36592 96988 36644
rect 97040 36632 97046 36644
rect 197446 36632 197452 36644
rect 97040 36604 197452 36632
rect 97040 36592 97046 36604
rect 197446 36592 197452 36604
rect 197504 36592 197510 36644
rect 118234 36524 118240 36576
rect 118292 36564 118298 36576
rect 408494 36564 408500 36576
rect 118292 36536 408500 36564
rect 118292 36524 118298 36536
rect 408494 36524 408500 36536
rect 408552 36524 408558 36576
rect 115198 35436 115204 35488
rect 115256 35476 115262 35488
rect 418154 35476 418160 35488
rect 115256 35448 418160 35476
rect 115256 35436 115262 35448
rect 418154 35436 418160 35448
rect 418212 35436 418218 35488
rect 117498 35368 117504 35420
rect 117556 35408 117562 35420
rect 440326 35408 440332 35420
rect 117556 35380 440332 35408
rect 117556 35368 117562 35380
rect 440326 35368 440332 35380
rect 440384 35368 440390 35420
rect 117406 35300 117412 35352
rect 117464 35340 117470 35352
rect 444374 35340 444380 35352
rect 117464 35312 444380 35340
rect 117464 35300 117470 35312
rect 444374 35300 444380 35312
rect 444432 35300 444438 35352
rect 120718 35232 120724 35284
rect 120776 35272 120782 35284
rect 478874 35272 478880 35284
rect 120776 35244 478880 35272
rect 120776 35232 120782 35244
rect 478874 35232 478880 35244
rect 478932 35232 478938 35284
rect 124858 35164 124864 35216
rect 124916 35204 124922 35216
rect 531314 35204 531320 35216
rect 124916 35176 531320 35204
rect 124916 35164 124922 35176
rect 531314 35164 531320 35176
rect 531372 35164 531378 35216
rect 111058 34280 111064 34332
rect 111116 34320 111122 34332
rect 363046 34320 363052 34332
rect 111116 34292 363052 34320
rect 111116 34280 111122 34292
rect 363046 34280 363052 34292
rect 363104 34280 363110 34332
rect 110966 34212 110972 34264
rect 111024 34252 111030 34264
rect 365714 34252 365720 34264
rect 111024 34224 365720 34252
rect 111024 34212 111030 34224
rect 365714 34212 365720 34224
rect 365772 34212 365778 34264
rect 115106 34144 115112 34196
rect 115164 34184 115170 34196
rect 407206 34184 407212 34196
rect 115164 34156 407212 34184
rect 115164 34144 115170 34156
rect 407206 34144 407212 34156
rect 407264 34144 407270 34196
rect 115014 34076 115020 34128
rect 115072 34116 115078 34128
rect 411254 34116 411260 34128
rect 115072 34088 411260 34116
rect 115072 34076 115078 34088
rect 411254 34076 411260 34088
rect 411312 34076 411318 34128
rect 114922 34008 114928 34060
rect 114980 34048 114986 34060
rect 414014 34048 414020 34060
rect 114980 34020 414020 34048
rect 114980 34008 114986 34020
rect 414014 34008 414020 34020
rect 414072 34008 414078 34060
rect 116026 33940 116032 33992
rect 116084 33980 116090 33992
rect 427814 33980 427820 33992
rect 116084 33952 427820 33980
rect 116084 33940 116090 33952
rect 427814 33940 427820 33952
rect 427872 33940 427878 33992
rect 116118 33872 116124 33924
rect 116176 33912 116182 33924
rect 430574 33912 430580 33924
rect 116176 33884 430580 33912
rect 116176 33872 116182 33884
rect 430574 33872 430580 33884
rect 430632 33872 430638 33924
rect 117314 33804 117320 33856
rect 117372 33844 117378 33856
rect 447134 33844 447140 33856
rect 117372 33816 447140 33844
rect 117372 33804 117378 33816
rect 447134 33804 447140 33816
rect 447192 33804 447198 33856
rect 120626 33736 120632 33788
rect 120684 33776 120690 33788
rect 481634 33776 481640 33788
rect 120684 33748 481640 33776
rect 120684 33736 120690 33748
rect 481634 33736 481640 33748
rect 481692 33736 481698 33788
rect 98362 32852 98368 32904
rect 98420 32892 98426 32904
rect 216674 32892 216680 32904
rect 98420 32864 216680 32892
rect 98420 32852 98426 32864
rect 216674 32852 216680 32864
rect 216732 32852 216738 32904
rect 108390 32784 108396 32836
rect 108448 32824 108454 32836
rect 332594 32824 332600 32836
rect 108448 32796 332600 32824
rect 108448 32784 108454 32796
rect 332594 32784 332600 32796
rect 332652 32784 332658 32836
rect 112254 32716 112260 32768
rect 112312 32756 112318 32768
rect 378134 32756 378140 32768
rect 112312 32728 378140 32756
rect 112312 32716 112318 32728
rect 378134 32716 378140 32728
rect 378192 32716 378198 32768
rect 112346 32648 112352 32700
rect 112404 32688 112410 32700
rect 380894 32688 380900 32700
rect 112404 32660 380900 32688
rect 112404 32648 112410 32660
rect 380894 32648 380900 32660
rect 380952 32648 380958 32700
rect 112162 32580 112168 32632
rect 112220 32620 112226 32632
rect 385126 32620 385132 32632
rect 112220 32592 385132 32620
rect 112220 32580 112226 32592
rect 385126 32580 385132 32592
rect 385184 32580 385190 32632
rect 113726 32512 113732 32564
rect 113784 32552 113790 32564
rect 390646 32552 390652 32564
rect 113784 32524 390652 32552
rect 113784 32512 113790 32524
rect 390646 32512 390652 32524
rect 390704 32512 390710 32564
rect 113634 32444 113640 32496
rect 113692 32484 113698 32496
rect 394694 32484 394700 32496
rect 113692 32456 394700 32484
rect 113692 32444 113698 32456
rect 394694 32444 394700 32456
rect 394752 32444 394758 32496
rect 113542 32376 113548 32428
rect 113600 32416 113606 32428
rect 397454 32416 397460 32428
rect 113600 32388 397460 32416
rect 113600 32376 113606 32388
rect 397454 32376 397460 32388
rect 397512 32376 397518 32428
rect 94038 31492 94044 31544
rect 94096 31532 94102 31544
rect 158806 31532 158812 31544
rect 94096 31504 158812 31532
rect 94096 31492 94102 31504
rect 158806 31492 158812 31504
rect 158864 31492 158870 31544
rect 94130 31424 94136 31476
rect 94188 31464 94194 31476
rect 162854 31464 162860 31476
rect 94188 31436 162860 31464
rect 94188 31424 94194 31436
rect 162854 31424 162860 31436
rect 162912 31424 162918 31476
rect 106918 31356 106924 31408
rect 106976 31396 106982 31408
rect 316034 31396 316040 31408
rect 106976 31368 316040 31396
rect 106976 31356 106982 31368
rect 316034 31356 316040 31368
rect 316092 31356 316098 31408
rect 108298 31288 108304 31340
rect 108356 31328 108362 31340
rect 325694 31328 325700 31340
rect 108356 31300 325700 31328
rect 108356 31288 108362 31300
rect 325694 31288 325700 31300
rect 325752 31288 325758 31340
rect 109494 31220 109500 31272
rect 109552 31260 109558 31272
rect 340966 31260 340972 31272
rect 109552 31232 340972 31260
rect 109552 31220 109558 31232
rect 340966 31220 340972 31232
rect 341024 31220 341030 31272
rect 111426 31152 111432 31204
rect 111484 31192 111490 31204
rect 354674 31192 354680 31204
rect 111484 31164 354680 31192
rect 111484 31152 111490 31164
rect 354674 31152 354680 31164
rect 354732 31152 354738 31204
rect 110782 31084 110788 31136
rect 110840 31124 110846 31136
rect 361574 31124 361580 31136
rect 110840 31096 361580 31124
rect 110840 31084 110846 31096
rect 361574 31084 361580 31096
rect 361632 31084 361638 31136
rect 110874 31016 110880 31068
rect 110932 31056 110938 31068
rect 364334 31056 364340 31068
rect 110932 31028 364340 31056
rect 110932 31016 110938 31028
rect 364334 31016 364340 31028
rect 364392 31016 364398 31068
rect 93946 30132 93952 30184
rect 94004 30172 94010 30184
rect 160094 30172 160100 30184
rect 94004 30144 160100 30172
rect 94004 30132 94010 30144
rect 160094 30132 160100 30144
rect 160152 30132 160158 30184
rect 106734 30064 106740 30116
rect 106792 30104 106798 30116
rect 307846 30104 307852 30116
rect 106792 30076 307852 30104
rect 106792 30064 106798 30076
rect 307846 30064 307852 30076
rect 307904 30064 307910 30116
rect 106826 29996 106832 30048
rect 106884 30036 106890 30048
rect 309134 30036 309140 30048
rect 106884 30008 309140 30036
rect 106884 29996 106890 30008
rect 309134 29996 309140 30008
rect 309192 29996 309198 30048
rect 106550 29928 106556 29980
rect 106608 29968 106614 29980
rect 311894 29968 311900 29980
rect 106608 29940 311900 29968
rect 106608 29928 106614 29940
rect 311894 29928 311900 29940
rect 311952 29928 311958 29980
rect 106642 29860 106648 29912
rect 106700 29900 106706 29912
rect 313366 29900 313372 29912
rect 106700 29872 313372 29900
rect 106700 29860 106706 29872
rect 313366 29860 313372 29872
rect 313424 29860 313430 29912
rect 106458 29792 106464 29844
rect 106516 29832 106522 29844
rect 314654 29832 314660 29844
rect 106516 29804 314660 29832
rect 106516 29792 106522 29804
rect 314654 29792 314660 29804
rect 314712 29792 314718 29844
rect 108114 29724 108120 29776
rect 108172 29764 108178 29776
rect 324406 29764 324412 29776
rect 108172 29736 324412 29764
rect 108172 29724 108178 29736
rect 324406 29724 324412 29736
rect 324464 29724 324470 29776
rect 108206 29656 108212 29708
rect 108264 29696 108270 29708
rect 328454 29696 328460 29708
rect 108264 29668 328460 29696
rect 108264 29656 108270 29668
rect 328454 29656 328460 29668
rect 328512 29656 328518 29708
rect 120534 29588 120540 29640
rect 120592 29628 120598 29640
rect 478966 29628 478972 29640
rect 120592 29600 478972 29628
rect 120592 29588 120598 29600
rect 478966 29588 478972 29600
rect 479024 29588 479030 29640
rect 104066 28636 104072 28688
rect 104124 28676 104130 28688
rect 276014 28676 276020 28688
rect 104124 28648 276020 28676
rect 104124 28636 104130 28648
rect 276014 28636 276020 28648
rect 276072 28636 276078 28688
rect 103974 28568 103980 28620
rect 104032 28608 104038 28620
rect 280154 28608 280160 28620
rect 104032 28580 280160 28608
rect 104032 28568 104038 28580
rect 280154 28568 280160 28580
rect 280212 28568 280218 28620
rect 104158 28500 104164 28552
rect 104216 28540 104222 28552
rect 281534 28540 281540 28552
rect 104216 28512 281540 28540
rect 104216 28500 104222 28512
rect 281534 28500 281540 28512
rect 281592 28500 281598 28552
rect 105354 28432 105360 28484
rect 105412 28472 105418 28484
rect 291286 28472 291292 28484
rect 105412 28444 291292 28472
rect 105412 28432 105418 28444
rect 291286 28432 291292 28444
rect 291344 28432 291350 28484
rect 105446 28364 105452 28416
rect 105504 28404 105510 28416
rect 295334 28404 295340 28416
rect 105504 28376 295340 28404
rect 105504 28364 105510 28376
rect 295334 28364 295340 28376
rect 295392 28364 295398 28416
rect 105262 28296 105268 28348
rect 105320 28336 105326 28348
rect 299474 28336 299480 28348
rect 105320 28308 299480 28336
rect 105320 28296 105326 28308
rect 299474 28296 299480 28308
rect 299532 28296 299538 28348
rect 110690 28228 110696 28280
rect 110748 28268 110754 28280
rect 357526 28268 357532 28280
rect 110748 28240 357532 28268
rect 110748 28228 110754 28240
rect 357526 28228 357532 28240
rect 357584 28228 357590 28280
rect 92842 27276 92848 27328
rect 92900 27316 92906 27328
rect 149054 27316 149060 27328
rect 92900 27288 149060 27316
rect 92900 27276 92906 27288
rect 149054 27276 149060 27288
rect 149112 27276 149118 27328
rect 92934 27208 92940 27260
rect 92992 27248 92998 27260
rect 150434 27248 150440 27260
rect 92992 27220 150440 27248
rect 92992 27208 92998 27220
rect 150434 27208 150440 27220
rect 150492 27208 150498 27260
rect 102870 27140 102876 27192
rect 102928 27180 102934 27192
rect 258166 27180 258172 27192
rect 102928 27152 258172 27180
rect 102928 27140 102934 27152
rect 258166 27140 258172 27152
rect 258224 27140 258230 27192
rect 102686 27072 102692 27124
rect 102744 27112 102750 27124
rect 262214 27112 262220 27124
rect 102744 27084 262220 27112
rect 102744 27072 102750 27084
rect 262214 27072 262220 27084
rect 262272 27072 262278 27124
rect 102778 27004 102784 27056
rect 102836 27044 102842 27056
rect 264974 27044 264980 27056
rect 102836 27016 264980 27044
rect 102836 27004 102842 27016
rect 264974 27004 264980 27016
rect 265032 27004 265038 27056
rect 103882 26936 103888 26988
rect 103940 26976 103946 26988
rect 274726 26976 274732 26988
rect 103940 26948 274732 26976
rect 103940 26936 103946 26948
rect 274726 26936 274732 26948
rect 274784 26936 274790 26988
rect 103790 26868 103796 26920
rect 103848 26908 103854 26920
rect 278774 26908 278780 26920
rect 103848 26880 278780 26908
rect 103848 26868 103854 26880
rect 278774 26868 278780 26880
rect 278832 26868 278838 26920
rect 92750 26052 92756 26104
rect 92808 26092 92814 26104
rect 146294 26092 146300 26104
rect 92808 26064 146300 26092
rect 92808 26052 92814 26064
rect 146294 26052 146300 26064
rect 146352 26052 146358 26104
rect 100846 25984 100852 26036
rect 100904 26024 100910 26036
rect 241606 26024 241612 26036
rect 100904 25996 241612 26024
rect 100904 25984 100910 25996
rect 241606 25984 241612 25996
rect 241664 25984 241670 26036
rect 101122 25916 101128 25968
rect 101180 25956 101186 25968
rect 245654 25956 245660 25968
rect 101180 25928 245660 25956
rect 101180 25916 101186 25928
rect 245654 25916 245660 25928
rect 245712 25916 245718 25968
rect 100938 25848 100944 25900
rect 100996 25888 101002 25900
rect 248414 25888 248420 25900
rect 100996 25860 248420 25888
rect 100996 25848 101002 25860
rect 248414 25848 248420 25860
rect 248472 25848 248478 25900
rect 101030 25780 101036 25832
rect 101088 25820 101094 25832
rect 252646 25820 252652 25832
rect 101088 25792 252652 25820
rect 101088 25780 101094 25792
rect 252646 25780 252652 25792
rect 252704 25780 252710 25832
rect 111886 25712 111892 25764
rect 111944 25752 111950 25764
rect 375374 25752 375380 25764
rect 111944 25724 375380 25752
rect 111944 25712 111950 25724
rect 375374 25712 375380 25724
rect 375432 25712 375438 25764
rect 111978 25644 111984 25696
rect 112036 25684 112042 25696
rect 379606 25684 379612 25696
rect 112036 25656 379612 25684
rect 112036 25644 112042 25656
rect 379606 25644 379612 25656
rect 379664 25644 379670 25696
rect 112070 25576 112076 25628
rect 112128 25616 112134 25628
rect 382274 25616 382280 25628
rect 112128 25588 382280 25616
rect 112128 25576 112134 25588
rect 382274 25576 382280 25588
rect 382332 25576 382338 25628
rect 113450 25508 113456 25560
rect 113508 25548 113514 25560
rect 396074 25548 396080 25560
rect 113508 25520 396080 25548
rect 113508 25508 113514 25520
rect 396074 25508 396080 25520
rect 396132 25508 396138 25560
rect 92658 24488 92664 24540
rect 92716 24528 92722 24540
rect 142246 24528 142252 24540
rect 92716 24500 142252 24528
rect 92716 24488 92722 24500
rect 142246 24488 142252 24500
rect 142304 24488 142310 24540
rect 96890 24420 96896 24472
rect 96948 24460 96954 24472
rect 198734 24460 198740 24472
rect 96948 24432 198740 24460
rect 96948 24420 96954 24432
rect 198734 24420 198740 24432
rect 198792 24420 198798 24472
rect 98178 24352 98184 24404
rect 98236 24392 98242 24404
rect 208486 24392 208492 24404
rect 98236 24364 208492 24392
rect 98236 24352 98242 24364
rect 208486 24352 208492 24364
rect 208544 24352 208550 24404
rect 98086 24284 98092 24336
rect 98144 24324 98150 24336
rect 212534 24324 212540 24336
rect 98144 24296 212540 24324
rect 98144 24284 98150 24296
rect 212534 24284 212540 24296
rect 212592 24284 212598 24336
rect 98270 24216 98276 24268
rect 98328 24256 98334 24268
rect 215294 24256 215300 24268
rect 98328 24228 215300 24256
rect 98328 24216 98334 24228
rect 215294 24216 215300 24228
rect 215352 24216 215358 24268
rect 110598 24148 110604 24200
rect 110656 24188 110662 24200
rect 358814 24188 358820 24200
rect 110656 24160 358820 24188
rect 110656 24148 110662 24160
rect 358814 24148 358820 24160
rect 358872 24148 358878 24200
rect 118970 24080 118976 24132
rect 119028 24120 119034 24132
rect 463694 24120 463700 24132
rect 119028 24092 463700 24120
rect 119028 24080 119034 24092
rect 463694 24080 463700 24092
rect 463752 24080 463758 24132
rect 95602 23128 95608 23180
rect 95660 23168 95666 23180
rect 179414 23168 179420 23180
rect 95660 23140 179420 23168
rect 95660 23128 95666 23140
rect 179414 23128 179420 23140
rect 179472 23128 179478 23180
rect 95510 23060 95516 23112
rect 95568 23100 95574 23112
rect 182174 23100 182180 23112
rect 95568 23072 182180 23100
rect 95568 23060 95574 23072
rect 182174 23060 182180 23072
rect 182232 23060 182238 23112
rect 96798 22992 96804 23044
rect 96856 23032 96862 23044
rect 191926 23032 191932 23044
rect 96856 23004 191932 23032
rect 96856 22992 96862 23004
rect 191926 22992 191932 23004
rect 191984 22992 191990 23044
rect 96706 22924 96712 22976
rect 96764 22964 96770 22976
rect 195974 22964 195980 22976
rect 96764 22936 195980 22964
rect 96764 22924 96770 22936
rect 195974 22924 195980 22936
rect 196032 22924 196038 22976
rect 100754 22856 100760 22908
rect 100812 22896 100818 22908
rect 249794 22896 249800 22908
rect 100812 22868 249800 22896
rect 100812 22856 100818 22868
rect 249794 22856 249800 22868
rect 249852 22856 249858 22908
rect 102594 22788 102600 22840
rect 102652 22828 102658 22840
rect 259454 22828 259460 22840
rect 102652 22800 259460 22828
rect 102652 22788 102658 22800
rect 259454 22788 259460 22800
rect 259512 22788 259518 22840
rect 102502 22720 102508 22772
rect 102560 22760 102566 22772
rect 263594 22760 263600 22772
rect 102560 22732 263600 22760
rect 102560 22720 102566 22732
rect 263594 22720 263600 22732
rect 263652 22720 263658 22772
rect 93578 21836 93584 21888
rect 93636 21876 93642 21888
rect 147674 21876 147680 21888
rect 93636 21848 147680 21876
rect 93636 21836 93642 21848
rect 147674 21836 147680 21848
rect 147732 21836 147738 21888
rect 95418 21768 95424 21820
rect 95476 21808 95482 21820
rect 175366 21808 175372 21820
rect 95476 21780 175372 21808
rect 95476 21768 95482 21780
rect 175366 21768 175372 21780
rect 175424 21768 175430 21820
rect 99558 21700 99564 21752
rect 99616 21740 99622 21752
rect 226334 21740 226340 21752
rect 99616 21712 226340 21740
rect 99616 21700 99622 21712
rect 226334 21700 226340 21712
rect 226392 21700 226398 21752
rect 123294 21632 123300 21684
rect 123352 21672 123358 21684
rect 506566 21672 506572 21684
rect 123352 21644 506572 21672
rect 123352 21632 123358 21644
rect 506566 21632 506572 21644
rect 506624 21632 506630 21684
rect 123202 21564 123208 21616
rect 123260 21604 123266 21616
rect 510614 21604 510620 21616
rect 123260 21576 510620 21604
rect 123260 21564 123266 21576
rect 510614 21564 510620 21576
rect 510672 21564 510678 21616
rect 123110 21496 123116 21548
rect 123168 21536 123174 21548
rect 513374 21536 513380 21548
rect 123168 21508 513380 21536
rect 123168 21496 123174 21508
rect 513374 21496 513380 21508
rect 513432 21496 513438 21548
rect 124766 21428 124772 21480
rect 124824 21468 124830 21480
rect 523126 21468 523132 21480
rect 124824 21440 523132 21468
rect 124824 21428 124830 21440
rect 523126 21428 523132 21440
rect 523184 21428 523190 21480
rect 38654 21360 38660 21412
rect 38712 21400 38718 21412
rect 83642 21400 83648 21412
rect 38712 21372 83648 21400
rect 38712 21360 38718 21372
rect 83642 21360 83648 21372
rect 83700 21360 83706 21412
rect 90266 21360 90272 21412
rect 90324 21400 90330 21412
rect 110598 21400 110604 21412
rect 90324 21372 110604 21400
rect 90324 21360 90330 21372
rect 110598 21360 110604 21372
rect 110656 21360 110662 21412
rect 126146 21360 126152 21412
rect 126204 21400 126210 21412
rect 550634 21400 550640 21412
rect 126204 21372 550640 21400
rect 126204 21360 126210 21372
rect 550634 21360 550640 21372
rect 550692 21360 550698 21412
rect 97994 20408 98000 20460
rect 98052 20448 98058 20460
rect 213914 20448 213920 20460
rect 98052 20420 213920 20448
rect 98052 20408 98058 20420
rect 213914 20408 213920 20420
rect 213972 20408 213978 20460
rect 122098 20340 122104 20392
rect 122156 20380 122162 20392
rect 490006 20380 490012 20392
rect 122156 20352 490012 20380
rect 122156 20340 122162 20352
rect 490006 20340 490012 20352
rect 490064 20340 490070 20392
rect 122006 20272 122012 20324
rect 122064 20312 122070 20324
rect 494054 20312 494060 20324
rect 122064 20284 494060 20312
rect 122064 20272 122070 20284
rect 494054 20272 494060 20284
rect 494112 20272 494118 20324
rect 122190 20204 122196 20256
rect 122248 20244 122254 20256
rect 496814 20244 496820 20256
rect 122248 20216 496820 20244
rect 122248 20204 122254 20216
rect 496814 20204 496820 20216
rect 496872 20204 496878 20256
rect 121914 20136 121920 20188
rect 121972 20176 121978 20188
rect 500954 20176 500960 20188
rect 121972 20148 500960 20176
rect 121972 20136 121978 20148
rect 500954 20136 500960 20148
rect 501012 20136 501018 20188
rect 126054 20068 126060 20120
rect 126112 20108 126118 20120
rect 546494 20108 546500 20120
rect 126112 20080 546500 20108
rect 126112 20068 126118 20080
rect 546494 20068 546500 20080
rect 546552 20068 546558 20120
rect 84746 20000 84752 20052
rect 84804 20040 84810 20052
rect 87782 20040 87788 20052
rect 84804 20012 87788 20040
rect 84804 20000 84810 20012
rect 87782 20000 87788 20012
rect 87840 20000 87846 20052
rect 127802 20000 127808 20052
rect 127860 20040 127866 20052
rect 557534 20040 557540 20052
rect 127860 20012 557540 20040
rect 127860 20000 127866 20012
rect 557534 20000 557540 20012
rect 557592 20000 557598 20052
rect 89070 19932 89076 19984
rect 89128 19972 89134 19984
rect 98086 19972 98092 19984
rect 89128 19944 98092 19972
rect 89128 19932 89134 19944
rect 98086 19932 98092 19944
rect 98144 19932 98150 19984
rect 127434 19932 127440 19984
rect 127492 19972 127498 19984
rect 561674 19972 561680 19984
rect 127492 19944 561680 19972
rect 127492 19932 127498 19944
rect 561674 19932 561680 19944
rect 561732 19932 561738 19984
rect 114830 18980 114836 19032
rect 114888 19020 114894 19032
rect 169018 19020 169024 19032
rect 114888 18992 169024 19020
rect 114888 18980 114894 18992
rect 169018 18980 169024 18992
rect 169076 18980 169082 19032
rect 93854 18912 93860 18964
rect 93912 18952 93918 18964
rect 168374 18952 168380 18964
rect 93912 18924 168380 18952
rect 93912 18912 93918 18924
rect 168374 18912 168380 18924
rect 168432 18912 168438 18964
rect 96338 18844 96344 18896
rect 96396 18884 96402 18896
rect 183554 18884 183560 18896
rect 96396 18856 183560 18884
rect 96396 18844 96402 18856
rect 183554 18844 183560 18856
rect 183612 18844 183618 18896
rect 118878 18776 118884 18828
rect 118936 18816 118942 18828
rect 466454 18816 466460 18828
rect 118936 18788 466460 18816
rect 118936 18776 118942 18788
rect 466454 18776 466460 18788
rect 466512 18776 466518 18828
rect 120442 18708 120448 18760
rect 120500 18748 120506 18760
rect 477494 18748 477500 18760
rect 120500 18720 477500 18748
rect 120500 18708 120506 18720
rect 477494 18708 477500 18720
rect 477552 18708 477558 18760
rect 123018 18640 123024 18692
rect 123076 18680 123082 18692
rect 517514 18680 517520 18692
rect 123076 18652 517520 18680
rect 123076 18640 123082 18652
rect 517514 18640 517520 18652
rect 517572 18640 517578 18692
rect 124674 18572 124680 18624
rect 124732 18612 124738 18624
rect 524414 18612 524420 18624
rect 124732 18584 524420 18612
rect 124732 18572 124738 18584
rect 524414 18572 524420 18584
rect 524472 18572 524478 18624
rect 93026 17620 93032 17672
rect 93084 17660 93090 17672
rect 143534 17660 143540 17672
rect 93084 17632 143540 17660
rect 93084 17620 93090 17632
rect 143534 17620 143540 17632
rect 143592 17620 143598 17672
rect 94682 17552 94688 17604
rect 94740 17592 94746 17604
rect 164326 17592 164332 17604
rect 94740 17564 164332 17592
rect 94740 17552 94746 17564
rect 164326 17552 164332 17564
rect 164384 17552 164390 17604
rect 118694 17484 118700 17536
rect 118752 17524 118758 17536
rect 459554 17524 459560 17536
rect 118752 17496 459560 17524
rect 118752 17484 118758 17496
rect 459554 17484 459560 17496
rect 459612 17484 459618 17536
rect 118786 17416 118792 17468
rect 118844 17456 118850 17468
rect 462406 17456 462412 17468
rect 118844 17428 462412 17456
rect 118844 17416 118850 17428
rect 462406 17416 462412 17428
rect 462464 17416 462470 17468
rect 120350 17348 120356 17400
rect 120408 17388 120414 17400
rect 474734 17388 474740 17400
rect 120408 17360 474740 17388
rect 120408 17348 120414 17360
rect 474734 17348 474740 17360
rect 474792 17348 474798 17400
rect 121822 17280 121828 17332
rect 121880 17320 121886 17332
rect 491294 17320 491300 17332
rect 121880 17292 491300 17320
rect 121880 17280 121886 17292
rect 491294 17280 491300 17292
rect 491352 17280 491358 17332
rect 121730 17212 121736 17264
rect 121788 17252 121794 17264
rect 495526 17252 495532 17264
rect 121788 17224 495532 17252
rect 121788 17212 121794 17224
rect 495526 17212 495532 17224
rect 495584 17212 495590 17264
rect 94590 16260 94596 16312
rect 94648 16300 94654 16312
rect 162026 16300 162032 16312
rect 94648 16272 162032 16300
rect 94648 16260 94654 16272
rect 162026 16260 162032 16272
rect 162084 16260 162090 16312
rect 114646 16192 114652 16244
rect 114704 16232 114710 16244
rect 412726 16232 412732 16244
rect 114704 16204 412732 16232
rect 114704 16192 114710 16204
rect 412726 16192 412732 16204
rect 412784 16192 412790 16244
rect 114738 16124 114744 16176
rect 114796 16164 114802 16176
rect 417234 16164 417240 16176
rect 114796 16136 417240 16164
rect 114796 16124 114802 16136
rect 417234 16124 417240 16136
rect 417292 16124 417298 16176
rect 114554 16056 114560 16108
rect 114612 16096 114618 16108
rect 418338 16096 418344 16108
rect 114612 16068 418344 16096
rect 114612 16056 114618 16068
rect 418338 16056 418344 16068
rect 418396 16056 418402 16108
rect 115934 15988 115940 16040
rect 115992 16028 115998 16040
rect 423766 16028 423772 16040
rect 115992 16000 423772 16028
rect 115992 15988 115998 16000
rect 423766 15988 423772 16000
rect 423824 15988 423830 16040
rect 125962 15920 125968 15972
rect 126020 15960 126026 15972
rect 541986 15960 541992 15972
rect 126020 15932 541992 15960
rect 126020 15920 126026 15932
rect 541986 15920 541992 15932
rect 542044 15920 542050 15972
rect 127710 15852 127716 15904
rect 127768 15892 127774 15904
rect 560754 15892 560760 15904
rect 127768 15864 560760 15892
rect 127768 15852 127774 15864
rect 560754 15852 560760 15864
rect 560812 15852 560818 15904
rect 109402 14764 109408 14816
rect 109460 14804 109466 14816
rect 352098 14804 352104 14816
rect 109460 14776 352104 14804
rect 109460 14764 109466 14776
rect 352098 14764 352104 14776
rect 352156 14764 352162 14816
rect 110506 14696 110512 14748
rect 110564 14736 110570 14748
rect 368658 14736 368664 14748
rect 110564 14708 368664 14736
rect 110564 14696 110570 14708
rect 368658 14696 368664 14708
rect 368716 14696 368722 14748
rect 111794 14628 111800 14680
rect 111852 14668 111858 14680
rect 384114 14668 384120 14680
rect 111852 14640 384120 14668
rect 111852 14628 111858 14640
rect 384114 14628 384120 14640
rect 384172 14628 384178 14680
rect 113358 14560 113364 14612
rect 113416 14600 113422 14612
rect 394050 14600 394056 14612
rect 113416 14572 394056 14600
rect 113416 14560 113422 14572
rect 394050 14560 394056 14572
rect 394108 14560 394114 14612
rect 113174 14492 113180 14544
rect 113232 14532 113238 14544
rect 396166 14532 396172 14544
rect 113232 14504 396172 14532
rect 113232 14492 113238 14504
rect 396166 14492 396172 14504
rect 396224 14492 396230 14544
rect 113266 14424 113272 14476
rect 113324 14464 113330 14476
rect 400674 14464 400680 14476
rect 113324 14436 400680 14464
rect 113324 14424 113330 14436
rect 400674 14424 400680 14436
rect 400732 14424 400738 14476
rect 93302 13472 93308 13524
rect 93360 13512 93366 13524
rect 155586 13512 155592 13524
rect 93360 13484 155592 13512
rect 93360 13472 93366 13484
rect 155586 13472 155592 13484
rect 155644 13472 155650 13524
rect 107930 13404 107936 13456
rect 107988 13444 107994 13456
rect 332226 13444 332232 13456
rect 107988 13416 332232 13444
rect 107988 13404 107994 13416
rect 332226 13404 332232 13416
rect 332284 13404 332290 13456
rect 108022 13336 108028 13388
rect 108080 13376 108086 13388
rect 335538 13376 335544 13388
rect 108080 13348 335544 13376
rect 108080 13336 108086 13348
rect 335538 13336 335544 13348
rect 335596 13336 335602 13388
rect 109126 13268 109132 13320
rect 109184 13308 109190 13320
rect 344370 13308 344376 13320
rect 109184 13280 344376 13308
rect 109184 13268 109190 13280
rect 344370 13268 344376 13280
rect 344428 13268 344434 13320
rect 109310 13200 109316 13252
rect 109368 13240 109374 13252
rect 346486 13240 346492 13252
rect 109368 13212 346492 13240
rect 109368 13200 109374 13212
rect 346486 13200 346492 13212
rect 346544 13200 346550 13252
rect 109218 13132 109224 13184
rect 109276 13172 109282 13184
rect 350994 13172 351000 13184
rect 109276 13144 351000 13172
rect 109276 13132 109282 13144
rect 350994 13132 351000 13144
rect 351052 13132 351058 13184
rect 110414 13064 110420 13116
rect 110472 13104 110478 13116
rect 367554 13104 367560 13116
rect 110472 13076 367560 13104
rect 110472 13064 110478 13076
rect 367554 13064 367560 13076
rect 367612 13064 367618 13116
rect 93210 12180 93216 12232
rect 93268 12220 93274 12232
rect 152274 12220 152280 12232
rect 93268 12192 152280 12220
rect 93268 12180 93274 12192
rect 152274 12180 152280 12192
rect 152332 12180 152338 12232
rect 106366 12112 106372 12164
rect 106424 12152 106430 12164
rect 317874 12152 317880 12164
rect 106424 12124 317880 12152
rect 106424 12112 106430 12124
rect 317874 12112 317880 12124
rect 317932 12112 317938 12164
rect 106274 12044 106280 12096
rect 106332 12084 106338 12096
rect 318978 12084 318984 12096
rect 106332 12056 318984 12084
rect 106332 12044 106338 12056
rect 318978 12044 318984 12056
rect 319036 12044 319042 12096
rect 107654 11976 107660 12028
rect 107712 12016 107718 12028
rect 327810 12016 327816 12028
rect 107712 11988 327816 12016
rect 107712 11976 107718 11988
rect 327810 11976 327816 11988
rect 327868 11976 327874 12028
rect 107838 11908 107844 11960
rect 107896 11948 107902 11960
rect 329926 11948 329932 11960
rect 107896 11920 329932 11948
rect 107896 11908 107902 11920
rect 329926 11908 329932 11920
rect 329984 11908 329990 11960
rect 107746 11840 107752 11892
rect 107804 11880 107810 11892
rect 334434 11880 334440 11892
rect 107804 11852 334440 11880
rect 107804 11840 107810 11852
rect 334434 11840 334440 11852
rect 334492 11840 334498 11892
rect 109034 11772 109040 11824
rect 109092 11812 109098 11824
rect 348786 11812 348792 11824
rect 109092 11784 348792 11812
rect 109092 11772 109098 11784
rect 348786 11772 348792 11784
rect 348844 11772 348850 11824
rect 125870 11704 125876 11756
rect 125928 11744 125934 11756
rect 544194 11744 544200 11756
rect 125928 11716 544200 11744
rect 125928 11704 125934 11716
rect 544194 11704 544200 11716
rect 544252 11704 544258 11756
rect 93118 10752 93124 10804
rect 93176 10792 93182 10804
rect 147766 10792 147772 10804
rect 93176 10764 147772 10792
rect 93176 10752 93182 10764
rect 147766 10752 147772 10764
rect 147824 10752 147830 10804
rect 102410 10684 102416 10736
rect 102468 10724 102474 10736
rect 269298 10724 269304 10736
rect 102468 10696 269304 10724
rect 102468 10684 102474 10696
rect 269298 10684 269304 10696
rect 269356 10684 269362 10736
rect 103698 10616 103704 10668
rect 103756 10656 103762 10668
rect 280246 10656 280252 10668
rect 103756 10628 280252 10656
rect 103756 10616 103762 10628
rect 280246 10616 280252 10628
rect 280304 10616 280310 10668
rect 103606 10548 103612 10600
rect 103664 10588 103670 10600
rect 284754 10588 284760 10600
rect 103664 10560 284760 10588
rect 103664 10548 103670 10560
rect 284754 10548 284760 10560
rect 284812 10548 284818 10600
rect 105078 10480 105084 10532
rect 105136 10520 105142 10532
rect 296806 10520 296812 10532
rect 105136 10492 296812 10520
rect 105136 10480 105142 10492
rect 296806 10480 296812 10492
rect 296864 10480 296870 10532
rect 104986 10412 104992 10464
rect 105044 10452 105050 10464
rect 301314 10452 301320 10464
rect 105044 10424 301320 10452
rect 105044 10412 105050 10424
rect 301314 10412 301320 10424
rect 301372 10412 301378 10464
rect 105170 10344 105176 10396
rect 105228 10384 105234 10396
rect 304626 10384 304632 10396
rect 105228 10356 304632 10384
rect 105228 10344 105234 10356
rect 304626 10344 304632 10356
rect 304684 10344 304690 10396
rect 125778 10276 125784 10328
rect 125836 10316 125842 10328
rect 539594 10316 539600 10328
rect 125836 10288 539600 10316
rect 125836 10276 125842 10288
rect 539594 10276 539600 10288
rect 539652 10276 539658 10328
rect 100570 9256 100576 9308
rect 100628 9296 100634 9308
rect 235074 9296 235080 9308
rect 100628 9268 235080 9296
rect 100628 9256 100634 9268
rect 235074 9256 235080 9268
rect 235132 9256 235138 9308
rect 102318 9188 102324 9240
rect 102376 9228 102382 9240
rect 261570 9228 261576 9240
rect 102376 9200 261576 9228
rect 102376 9188 102382 9200
rect 261570 9188 261576 9200
rect 261628 9188 261634 9240
rect 102134 9120 102140 9172
rect 102192 9160 102198 9172
rect 264882 9160 264888 9172
rect 102192 9132 264888 9160
rect 102192 9120 102198 9132
rect 264882 9120 264888 9132
rect 264940 9120 264946 9172
rect 102226 9052 102232 9104
rect 102284 9092 102290 9104
rect 268194 9092 268200 9104
rect 102284 9064 268200 9092
rect 102284 9052 102290 9064
rect 268194 9052 268200 9064
rect 268252 9052 268258 9104
rect 103514 8984 103520 9036
rect 103572 9024 103578 9036
rect 278130 9024 278136 9036
rect 103572 8996 278136 9024
rect 103572 8984 103578 8996
rect 278130 8984 278136 8996
rect 278188 8984 278194 9036
rect 209038 8916 209044 8968
rect 209096 8956 209102 8968
rect 557442 8956 557448 8968
rect 209096 8928 557448 8956
rect 209096 8916 209102 8928
rect 557442 8916 557448 8928
rect 557500 8916 557506 8968
rect 97534 8100 97540 8152
rect 97592 8140 97598 8152
rect 201954 8140 201960 8152
rect 97592 8112 201960 8140
rect 97592 8100 97598 8112
rect 201954 8100 201960 8112
rect 202012 8100 202018 8152
rect 96614 8032 96620 8084
rect 96672 8072 96678 8084
rect 205266 8072 205272 8084
rect 96672 8044 205272 8072
rect 96672 8032 96678 8044
rect 205266 8032 205272 8044
rect 205324 8032 205330 8084
rect 98822 7964 98828 8016
rect 98880 8004 98886 8016
rect 215202 8004 215208 8016
rect 98880 7976 215208 8004
rect 98880 7964 98886 7976
rect 215202 7964 215208 7976
rect 215260 7964 215266 8016
rect 99282 7896 99288 7948
rect 99340 7936 99346 7948
rect 221826 7936 221832 7948
rect 99340 7908 221832 7936
rect 99340 7896 99346 7908
rect 221826 7896 221832 7908
rect 221884 7896 221890 7948
rect 99466 7828 99472 7880
rect 99524 7868 99530 7880
rect 229554 7868 229560 7880
rect 99524 7840 229560 7868
rect 99524 7828 99530 7840
rect 229554 7828 229560 7840
rect 229612 7828 229618 7880
rect 100662 7760 100668 7812
rect 100720 7800 100726 7812
rect 231762 7800 231768 7812
rect 100720 7772 231768 7800
rect 100720 7760 100726 7772
rect 231762 7760 231768 7772
rect 231820 7760 231826 7812
rect 124582 7692 124588 7744
rect 124640 7732 124646 7744
rect 527634 7732 527640 7744
rect 124640 7704 527640 7732
rect 124640 7692 124646 7704
rect 527634 7692 527640 7704
rect 527692 7692 527698 7744
rect 61746 7624 61752 7676
rect 61804 7664 61810 7676
rect 86310 7664 86316 7676
rect 61804 7636 86316 7664
rect 61804 7624 61810 7636
rect 86310 7624 86316 7636
rect 86368 7624 86374 7676
rect 124490 7624 124496 7676
rect 124548 7664 124554 7676
rect 530946 7664 530952 7676
rect 124548 7636 530952 7664
rect 124548 7624 124554 7636
rect 530946 7624 530952 7636
rect 531004 7624 531010 7676
rect 26418 7556 26424 7608
rect 26476 7596 26482 7608
rect 83458 7596 83464 7608
rect 26476 7568 83464 7596
rect 26476 7556 26482 7568
rect 83458 7556 83464 7568
rect 83516 7556 83522 7608
rect 124398 7556 124404 7608
rect 124456 7596 124462 7608
rect 534258 7596 534264 7608
rect 124456 7568 534264 7596
rect 124456 7556 124462 7568
rect 534258 7556 534264 7568
rect 534316 7556 534322 7608
rect 517514 7488 517520 7540
rect 517572 7528 517578 7540
rect 518802 7528 518808 7540
rect 517572 7500 518808 7528
rect 517572 7488 517578 7500
rect 518802 7488 518808 7500
rect 518860 7488 518866 7540
rect 523126 7488 523132 7540
rect 523184 7528 523190 7540
rect 524322 7528 524328 7540
rect 523184 7500 524328 7528
rect 523184 7488 523190 7500
rect 524322 7488 524328 7500
rect 524380 7488 524386 7540
rect 73890 6740 73896 6792
rect 73948 6780 73954 6792
rect 85942 6780 85948 6792
rect 73948 6752 85948 6780
rect 73948 6740 73954 6752
rect 85942 6740 85948 6752
rect 86000 6740 86006 6792
rect 70578 6672 70584 6724
rect 70636 6712 70642 6724
rect 84930 6712 84936 6724
rect 70636 6684 84936 6712
rect 70636 6672 70642 6684
rect 84930 6672 84936 6684
rect 84988 6672 84994 6724
rect 68370 6604 68376 6656
rect 68428 6644 68434 6656
rect 86034 6644 86040 6656
rect 68428 6616 86040 6644
rect 68428 6604 68434 6616
rect 86034 6604 86040 6616
rect 86092 6604 86098 6656
rect 67266 6536 67272 6588
rect 67324 6576 67330 6588
rect 86218 6576 86224 6588
rect 67324 6548 86224 6576
rect 67324 6536 67330 6548
rect 86218 6536 86224 6548
rect 86276 6536 86282 6588
rect 91186 6536 91192 6588
rect 91244 6576 91250 6588
rect 129090 6576 129096 6588
rect 91244 6548 129096 6576
rect 91244 6536 91250 6548
rect 129090 6536 129096 6548
rect 129148 6536 129154 6588
rect 63954 6468 63960 6520
rect 64012 6508 64018 6520
rect 86126 6508 86132 6520
rect 64012 6480 86132 6508
rect 64012 6468 64018 6480
rect 86126 6468 86132 6480
rect 86184 6468 86190 6520
rect 96062 6468 96068 6520
rect 96120 6508 96126 6520
rect 185394 6508 185400 6520
rect 96120 6480 185400 6508
rect 96120 6468 96126 6480
rect 185394 6468 185400 6480
rect 185452 6468 185458 6520
rect 62850 6400 62856 6452
rect 62908 6440 62914 6452
rect 84838 6440 84844 6452
rect 62908 6412 84844 6440
rect 62908 6400 62914 6412
rect 84838 6400 84844 6412
rect 84896 6400 84902 6452
rect 95970 6400 95976 6452
rect 96028 6440 96034 6452
rect 188706 6440 188712 6452
rect 96028 6412 188712 6440
rect 96028 6400 96034 6412
rect 188706 6400 188712 6412
rect 188764 6400 188770 6452
rect 55122 6332 55128 6384
rect 55180 6372 55186 6384
rect 84654 6372 84660 6384
rect 55180 6344 84660 6372
rect 55180 6332 55186 6344
rect 84654 6332 84660 6344
rect 84712 6332 84718 6384
rect 91830 6332 91836 6384
rect 91888 6372 91894 6384
rect 106182 6372 106188 6384
rect 91888 6344 106188 6372
rect 91888 6332 91894 6344
rect 106182 6332 106188 6344
rect 106240 6332 106246 6384
rect 122926 6332 122932 6384
rect 122984 6372 122990 6384
rect 517698 6372 517704 6384
rect 122984 6344 517704 6372
rect 122984 6332 122990 6344
rect 517698 6332 517704 6344
rect 517756 6332 517762 6384
rect 48498 6264 48504 6316
rect 48556 6304 48562 6316
rect 84562 6304 84568 6316
rect 48556 6276 84568 6304
rect 48556 6264 48562 6276
rect 84562 6264 84568 6276
rect 84620 6264 84626 6316
rect 91738 6264 91744 6316
rect 91796 6304 91802 6316
rect 114738 6304 114744 6316
rect 91796 6276 114744 6304
rect 91796 6264 91802 6276
rect 114738 6264 114744 6276
rect 114796 6264 114802 6316
rect 125686 6264 125692 6316
rect 125744 6304 125750 6316
rect 539778 6304 539784 6316
rect 125744 6276 539784 6304
rect 125744 6264 125750 6276
rect 539778 6264 539784 6276
rect 539836 6264 539842 6316
rect 38562 6196 38568 6248
rect 38620 6236 38626 6248
rect 83366 6236 83372 6248
rect 38620 6208 83372 6236
rect 38620 6196 38626 6208
rect 83366 6196 83372 6208
rect 83424 6196 83430 6248
rect 90174 6196 90180 6248
rect 90232 6236 90238 6248
rect 113634 6236 113640 6248
rect 90232 6208 113640 6236
rect 90232 6196 90238 6208
rect 113634 6196 113640 6208
rect 113692 6196 113698 6248
rect 127618 6196 127624 6248
rect 127676 6236 127682 6248
rect 556338 6236 556344 6248
rect 127676 6208 556344 6236
rect 127676 6196 127682 6208
rect 556338 6196 556344 6208
rect 556396 6196 556402 6248
rect 34146 6128 34152 6180
rect 34204 6168 34210 6180
rect 83274 6168 83280 6180
rect 34204 6140 83280 6168
rect 34204 6128 34210 6140
rect 83274 6128 83280 6140
rect 83332 6128 83338 6180
rect 90082 6128 90088 6180
rect 90140 6168 90146 6180
rect 116946 6168 116952 6180
rect 90140 6140 116952 6168
rect 90140 6128 90146 6140
rect 116946 6128 116952 6140
rect 117004 6128 117010 6180
rect 127526 6128 127532 6180
rect 127584 6168 127590 6180
rect 559650 6168 559656 6180
rect 127584 6140 559656 6168
rect 127584 6128 127590 6140
rect 559650 6128 559656 6140
rect 559708 6128 559714 6180
rect 88978 5448 88984 5500
rect 89036 5488 89042 5500
rect 100386 5488 100392 5500
rect 89036 5460 100392 5488
rect 89036 5448 89042 5460
rect 100386 5448 100392 5460
rect 100444 5448 100450 5500
rect 96246 5380 96252 5432
rect 96304 5420 96310 5432
rect 96304 5392 103514 5420
rect 96304 5380 96310 5392
rect 74994 5312 75000 5364
rect 75052 5352 75058 5364
rect 85850 5352 85856 5364
rect 75052 5324 85856 5352
rect 75052 5312 75058 5324
rect 85850 5312 85856 5324
rect 85908 5312 85914 5364
rect 90818 5312 90824 5364
rect 90876 5352 90882 5364
rect 103486 5352 103514 5392
rect 186498 5352 186504 5364
rect 90876 5324 98868 5352
rect 103486 5324 186504 5352
rect 90876 5312 90882 5324
rect 80054 5244 80060 5296
rect 80112 5284 80118 5296
rect 83182 5284 83188 5296
rect 80112 5256 83188 5284
rect 80112 5244 80118 5256
rect 83182 5244 83188 5256
rect 83240 5244 83246 5296
rect 88886 5244 88892 5296
rect 88944 5284 88950 5296
rect 97074 5284 97080 5296
rect 88944 5256 97080 5284
rect 88944 5244 88950 5256
rect 97074 5244 97080 5256
rect 97132 5244 97138 5296
rect 56226 5176 56232 5228
rect 56284 5216 56290 5228
rect 85022 5216 85028 5228
rect 56284 5188 85028 5216
rect 56284 5176 56290 5188
rect 85022 5176 85028 5188
rect 85080 5176 85086 5228
rect 89714 5176 89720 5228
rect 89772 5216 89778 5228
rect 98840 5216 98868 5324
rect 186498 5312 186504 5324
rect 186556 5312 186562 5364
rect 100110 5244 100116 5296
rect 100168 5284 100174 5296
rect 232866 5284 232872 5296
rect 100168 5256 232872 5284
rect 100168 5244 100174 5256
rect 232866 5244 232872 5256
rect 232924 5244 232930 5296
rect 103698 5216 103704 5228
rect 89772 5188 98684 5216
rect 98840 5188 103704 5216
rect 89772 5176 89778 5188
rect 52914 5108 52920 5160
rect 52972 5148 52978 5160
rect 85390 5148 85396 5160
rect 52972 5120 85396 5148
rect 52972 5108 52978 5120
rect 85390 5108 85396 5120
rect 85448 5108 85454 5160
rect 90450 5108 90456 5160
rect 90508 5148 90514 5160
rect 98656 5148 98684 5188
rect 103698 5176 103704 5188
rect 103756 5176 103762 5228
rect 104894 5176 104900 5228
rect 104952 5216 104958 5228
rect 299106 5216 299112 5228
rect 104952 5188 299112 5216
rect 104952 5176 104958 5188
rect 299106 5176 299112 5188
rect 299164 5176 299170 5228
rect 90508 5120 95832 5148
rect 98656 5120 98776 5148
rect 90508 5108 90514 5120
rect 50706 5040 50712 5092
rect 50764 5080 50770 5092
rect 85114 5080 85120 5092
rect 50764 5052 85120 5080
rect 50764 5040 50770 5052
rect 85114 5040 85120 5052
rect 85172 5040 85178 5092
rect 89990 5040 89996 5092
rect 90048 5080 90054 5092
rect 95804 5080 95832 5120
rect 98748 5080 98776 5120
rect 120166 5108 120172 5160
rect 120224 5148 120230 5160
rect 481266 5148 481272 5160
rect 120224 5120 481272 5148
rect 120224 5108 120230 5120
rect 481266 5108 481272 5120
rect 481324 5108 481330 5160
rect 107010 5080 107016 5092
rect 90048 5052 95648 5080
rect 95804 5052 98684 5080
rect 98748 5052 107016 5080
rect 90048 5040 90054 5052
rect 49602 4972 49608 5024
rect 49660 5012 49666 5024
rect 84470 5012 84476 5024
rect 49660 4984 84476 5012
rect 49660 4972 49666 4984
rect 84470 4972 84476 4984
rect 84528 4972 84534 5024
rect 25314 4904 25320 4956
rect 25372 4944 25378 4956
rect 82446 4944 82452 4956
rect 25372 4916 82452 4944
rect 25372 4904 25378 4916
rect 82446 4904 82452 4916
rect 82504 4904 82510 4956
rect 95620 4944 95648 5052
rect 98656 5012 98684 5052
rect 107010 5040 107016 5052
rect 107068 5040 107074 5092
rect 121638 5040 121644 5092
rect 121696 5080 121702 5092
rect 500034 5080 500040 5092
rect 121696 5052 500040 5080
rect 121696 5040 121702 5052
rect 500034 5040 500040 5052
rect 500092 5040 500098 5092
rect 108114 5012 108120 5024
rect 98656 4984 108120 5012
rect 108114 4972 108120 4984
rect 108172 4972 108178 5024
rect 122834 4972 122840 5024
rect 122892 5012 122898 5024
rect 509970 5012 509976 5024
rect 122892 4984 509976 5012
rect 122892 4972 122898 4984
rect 509970 4972 509976 4984
rect 510028 4972 510034 5024
rect 110322 4944 110328 4956
rect 95620 4916 110328 4944
rect 110322 4904 110328 4916
rect 110380 4904 110386 4956
rect 124306 4904 124312 4956
rect 124364 4944 124370 4956
rect 526530 4944 526536 4956
rect 124364 4916 526536 4944
rect 124364 4904 124370 4916
rect 526530 4904 526536 4916
rect 526588 4904 526594 4956
rect 24210 4836 24216 4888
rect 24268 4876 24274 4888
rect 81618 4876 81624 4888
rect 24268 4848 81624 4876
rect 24268 4836 24274 4848
rect 81618 4836 81624 4848
rect 81676 4836 81682 4888
rect 92014 4836 92020 4888
rect 92072 4876 92078 4888
rect 119154 4876 119160 4888
rect 92072 4848 119160 4876
rect 92072 4836 92078 4848
rect 119154 4836 119160 4848
rect 119212 4836 119218 4888
rect 124214 4836 124220 4888
rect 124272 4876 124278 4888
rect 516778 4876 516784 4888
rect 124272 4848 516784 4876
rect 124272 4836 124278 4848
rect 516778 4836 516784 4848
rect 516836 4836 516842 4888
rect 516888 4848 521654 4876
rect 23106 4768 23112 4820
rect 23164 4808 23170 4820
rect 81526 4808 81532 4820
rect 23164 4780 81532 4808
rect 23164 4768 23170 4780
rect 81526 4768 81532 4780
rect 81584 4768 81590 4820
rect 82354 4768 82360 4820
rect 82412 4808 82418 4820
rect 87690 4808 87696 4820
rect 82412 4780 87696 4808
rect 82412 4768 82418 4780
rect 87690 4768 87696 4780
rect 87748 4768 87754 4820
rect 89898 4768 89904 4820
rect 89956 4808 89962 4820
rect 120258 4808 120264 4820
rect 89956 4780 120264 4808
rect 89956 4768 89962 4780
rect 120258 4768 120264 4780
rect 120316 4768 120322 4820
rect 125594 4768 125600 4820
rect 125652 4808 125658 4820
rect 516888 4808 516916 4848
rect 125652 4780 516916 4808
rect 521626 4808 521654 4848
rect 548610 4808 548616 4820
rect 521626 4780 548616 4808
rect 125652 4768 125658 4780
rect 548610 4768 548616 4780
rect 548668 4768 548674 4820
rect 516778 4700 516784 4752
rect 516836 4740 516842 4752
rect 529842 4740 529848 4752
rect 516836 4712 529848 4740
rect 516836 4700 516842 4712
rect 529842 4700 529848 4712
rect 529900 4700 529906 4752
rect 88702 4292 88708 4344
rect 88760 4332 88766 4344
rect 94866 4332 94872 4344
rect 88760 4304 94872 4332
rect 88760 4292 88766 4304
rect 94866 4292 94872 4304
rect 94924 4292 94930 4344
rect 88794 4156 88800 4208
rect 88852 4196 88858 4208
rect 93762 4196 93768 4208
rect 88852 4168 93768 4196
rect 88852 4156 88858 4168
rect 93762 4156 93768 4168
rect 93820 4156 93826 4208
rect 75730 4088 75736 4140
rect 75788 4128 75794 4140
rect 83734 4128 83740 4140
rect 75788 4100 83740 4128
rect 75788 4088 75794 4100
rect 83734 4088 83740 4100
rect 83792 4088 83798 4140
rect 88426 4088 88432 4140
rect 88484 4128 88490 4140
rect 95970 4128 95976 4140
rect 88484 4100 95976 4128
rect 88484 4088 88490 4100
rect 95970 4088 95976 4100
rect 96028 4088 96034 4140
rect 131206 4088 131212 4140
rect 131264 4128 131270 4140
rect 132402 4128 132408 4140
rect 131264 4100 132408 4128
rect 131264 4088 131270 4100
rect 132402 4088 132408 4100
rect 132460 4088 132466 4140
rect 162118 4088 162124 4140
rect 162176 4128 162182 4140
rect 162176 4100 171134 4128
rect 162176 4088 162182 4100
rect 79410 4020 79416 4072
rect 79468 4060 79474 4072
rect 87506 4060 87512 4072
rect 79468 4032 87512 4060
rect 79468 4020 79474 4032
rect 87506 4020 87512 4032
rect 87564 4020 87570 4072
rect 98638 4020 98644 4072
rect 98696 4060 98702 4072
rect 170950 4060 170956 4072
rect 98696 4032 170956 4060
rect 98696 4020 98702 4032
rect 170950 4020 170956 4032
rect 171008 4020 171014 4072
rect 51810 3952 51816 4004
rect 51868 3992 51874 4004
rect 62758 3992 62764 4004
rect 51868 3964 62764 3992
rect 51868 3952 51874 3964
rect 62758 3952 62764 3964
rect 62816 3952 62822 4004
rect 76098 3952 76104 4004
rect 76156 3992 76162 4004
rect 87598 3992 87604 4004
rect 76156 3964 87604 3992
rect 76156 3952 76162 3964
rect 87598 3952 87604 3964
rect 87656 3952 87662 4004
rect 106182 3952 106188 4004
rect 106240 3992 106246 4004
rect 139026 3992 139032 4004
rect 106240 3964 139032 3992
rect 106240 3952 106246 3964
rect 139026 3952 139032 3964
rect 139084 3952 139090 4004
rect 142246 3952 142252 4004
rect 142304 3992 142310 4004
rect 143442 3992 143448 4004
rect 142304 3964 143448 3992
rect 142304 3952 142310 3964
rect 143442 3952 143448 3964
rect 143500 3952 143506 4004
rect 147766 3952 147772 4004
rect 147824 3992 147830 4004
rect 148962 3992 148968 4004
rect 147824 3964 148968 3992
rect 147824 3952 147830 3964
rect 148962 3952 148968 3964
rect 149020 3952 149026 4004
rect 158806 3952 158812 4004
rect 158864 3992 158870 4004
rect 160002 3992 160008 4004
rect 158864 3964 160008 3992
rect 158864 3952 158870 3964
rect 160002 3952 160008 3964
rect 160060 3952 160066 4004
rect 171106 3992 171134 4100
rect 175366 4020 175372 4072
rect 175424 4060 175430 4072
rect 176562 4060 176568 4072
rect 175424 4032 176568 4060
rect 175424 4020 175430 4032
rect 176562 4020 176568 4032
rect 176620 4020 176626 4072
rect 191926 4020 191932 4072
rect 191984 4060 191990 4072
rect 193122 4060 193128 4072
rect 191984 4032 193128 4060
rect 191984 4020 191990 4032
rect 193122 4020 193128 4032
rect 193180 4020 193186 4072
rect 208486 4020 208492 4072
rect 208544 4060 208550 4072
rect 209682 4060 209688 4072
rect 208544 4032 209688 4060
rect 208544 4020 208550 4032
rect 209682 4020 209688 4032
rect 209740 4020 209746 4072
rect 293586 4060 293592 4072
rect 277366 4032 293592 4060
rect 277366 3992 277394 4032
rect 293586 4020 293592 4032
rect 293644 4020 293650 4072
rect 296806 4020 296812 4072
rect 296864 4060 296870 4072
rect 298002 4060 298008 4072
rect 296864 4032 298008 4060
rect 296864 4020 296870 4032
rect 298002 4020 298008 4032
rect 298060 4020 298066 4072
rect 307846 4020 307852 4072
rect 307904 4060 307910 4072
rect 309042 4060 309048 4072
rect 307904 4032 309048 4060
rect 307904 4020 307910 4032
rect 309042 4020 309048 4032
rect 309100 4020 309106 4072
rect 324406 4020 324412 4072
rect 324464 4060 324470 4072
rect 325602 4060 325608 4072
rect 324464 4032 325608 4060
rect 324464 4020 324470 4032
rect 325602 4020 325608 4032
rect 325660 4020 325666 4072
rect 329926 4020 329932 4072
rect 329984 4060 329990 4072
rect 331122 4060 331128 4072
rect 329984 4032 331128 4060
rect 329984 4020 329990 4032
rect 331122 4020 331128 4032
rect 331180 4020 331186 4072
rect 340966 4020 340972 4072
rect 341024 4060 341030 4072
rect 342162 4060 342168 4072
rect 341024 4032 342168 4060
rect 341024 4020 341030 4032
rect 342162 4020 342168 4032
rect 342220 4020 342226 4072
rect 346486 4020 346492 4072
rect 346544 4060 346550 4072
rect 347682 4060 347688 4072
rect 346544 4032 347688 4060
rect 346544 4020 346550 4032
rect 347682 4020 347688 4032
rect 347740 4020 347746 4072
rect 357526 4020 357532 4072
rect 357584 4060 357590 4072
rect 358722 4060 358728 4072
rect 357584 4032 358728 4060
rect 357584 4020 357590 4032
rect 358722 4020 358728 4032
rect 358780 4020 358786 4072
rect 390646 4020 390652 4072
rect 390704 4060 390710 4072
rect 391842 4060 391848 4072
rect 390704 4032 391848 4060
rect 390704 4020 390710 4032
rect 391842 4020 391848 4032
rect 391900 4020 391906 4072
rect 396166 4020 396172 4072
rect 396224 4060 396230 4072
rect 397362 4060 397368 4072
rect 396224 4032 397368 4060
rect 396224 4020 396230 4032
rect 397362 4020 397368 4032
rect 397420 4020 397426 4072
rect 407206 4020 407212 4072
rect 407264 4060 407270 4072
rect 408402 4060 408408 4072
rect 407264 4032 408408 4060
rect 407264 4020 407270 4032
rect 408402 4020 408408 4032
rect 408460 4020 408466 4072
rect 161446 3964 164372 3992
rect 171106 3964 277394 3992
rect 44082 3884 44088 3936
rect 44140 3924 44146 3936
rect 54478 3924 54484 3936
rect 44140 3896 54484 3924
rect 44140 3884 44146 3896
rect 54478 3884 54484 3896
rect 54536 3884 54542 3936
rect 58434 3884 58440 3936
rect 58492 3924 58498 3936
rect 71038 3924 71044 3936
rect 58492 3896 71044 3924
rect 58492 3884 58498 3896
rect 71038 3884 71044 3896
rect 71096 3884 71102 3936
rect 72786 3884 72792 3936
rect 72844 3924 72850 3936
rect 86678 3924 86684 3936
rect 72844 3896 86684 3924
rect 72844 3884 72850 3896
rect 86678 3884 86684 3896
rect 86736 3884 86742 3936
rect 94498 3884 94504 3936
rect 94556 3924 94562 3936
rect 104802 3924 104808 3936
rect 94556 3896 104808 3924
rect 94556 3884 94562 3896
rect 104802 3884 104808 3896
rect 104860 3884 104866 3936
rect 115382 3884 115388 3936
rect 115440 3924 115446 3936
rect 135714 3924 135720 3936
rect 115440 3896 135720 3924
rect 115440 3884 115446 3896
rect 135714 3884 135720 3896
rect 135772 3884 135778 3936
rect 135990 3884 135996 3936
rect 136048 3924 136054 3936
rect 161446 3924 161474 3964
rect 136048 3896 161474 3924
rect 164344 3924 164372 3964
rect 278038 3952 278044 4004
rect 278096 3992 278102 4004
rect 278096 3964 287054 3992
rect 278096 3952 278102 3964
rect 210786 3924 210792 3936
rect 164344 3896 210792 3924
rect 136048 3884 136054 3896
rect 210786 3884 210792 3896
rect 210844 3884 210850 3936
rect 219526 3884 219532 3936
rect 219584 3924 219590 3936
rect 220722 3924 220728 3936
rect 219584 3896 220728 3924
rect 219584 3884 219590 3896
rect 220722 3884 220728 3896
rect 220780 3884 220786 3936
rect 225046 3884 225052 3936
rect 225104 3924 225110 3936
rect 226242 3924 226248 3936
rect 225104 3896 226248 3924
rect 225104 3884 225110 3896
rect 226242 3884 226248 3896
rect 226300 3884 226306 3936
rect 241606 3884 241612 3936
rect 241664 3924 241670 3936
rect 242802 3924 242808 3936
rect 241664 3896 242808 3924
rect 241664 3884 241670 3896
rect 242802 3884 242808 3896
rect 242860 3884 242866 3936
rect 247126 3884 247132 3936
rect 247184 3924 247190 3936
rect 248322 3924 248328 3936
rect 247184 3896 248328 3924
rect 247184 3884 247190 3896
rect 248322 3884 248328 3896
rect 248380 3884 248386 3936
rect 258166 3884 258172 3936
rect 258224 3924 258230 3936
rect 259362 3924 259368 3936
rect 258224 3896 259368 3924
rect 258224 3884 258230 3896
rect 259362 3884 259368 3896
rect 259420 3884 259426 3936
rect 274726 3884 274732 3936
rect 274784 3924 274790 3936
rect 275922 3924 275928 3936
rect 274784 3896 275928 3924
rect 274784 3884 274790 3896
rect 275922 3884 275928 3896
rect 275980 3884 275986 3936
rect 280246 3884 280252 3936
rect 280304 3924 280310 3936
rect 281442 3924 281448 3936
rect 280304 3896 281448 3924
rect 280304 3884 280310 3896
rect 281442 3884 281448 3896
rect 281500 3884 281506 3936
rect 287026 3924 287054 3964
rect 291286 3952 291292 4004
rect 291344 3992 291350 4004
rect 292482 3992 292488 4004
rect 291344 3964 292488 3992
rect 291344 3952 291350 3964
rect 292482 3952 292488 3964
rect 292540 3952 292546 4004
rect 295978 3952 295984 4004
rect 296036 3992 296042 4004
rect 469122 3992 469128 4004
rect 296036 3964 469128 3992
rect 296036 3952 296042 3964
rect 469122 3952 469128 3964
rect 469180 3952 469186 4004
rect 490098 3924 490104 3936
rect 287026 3896 490104 3924
rect 490098 3884 490104 3896
rect 490156 3884 490162 3936
rect 45186 3816 45192 3868
rect 45244 3856 45250 3868
rect 58618 3856 58624 3868
rect 45244 3828 58624 3856
rect 45244 3816 45250 3828
rect 58618 3816 58624 3828
rect 58676 3816 58682 3868
rect 69474 3816 69480 3868
rect 69532 3856 69538 3868
rect 86586 3856 86592 3868
rect 69532 3828 86592 3856
rect 69532 3816 69538 3828
rect 86586 3816 86592 3828
rect 86644 3816 86650 3868
rect 88334 3816 88340 3868
rect 88392 3856 88398 3868
rect 99282 3856 99288 3868
rect 88392 3828 99288 3856
rect 88392 3816 88398 3828
rect 99282 3816 99288 3828
rect 99340 3816 99346 3868
rect 128998 3816 129004 3868
rect 129056 3856 129062 3868
rect 164142 3856 164148 3868
rect 129056 3828 164148 3856
rect 129056 3816 129062 3828
rect 164142 3816 164148 3828
rect 164200 3816 164206 3868
rect 164326 3816 164332 3868
rect 164384 3856 164390 3868
rect 165522 3856 165528 3868
rect 164384 3828 165528 3856
rect 164384 3816 164390 3828
rect 165522 3816 165528 3828
rect 165580 3816 165586 3868
rect 169018 3816 169024 3868
rect 169076 3856 169082 3868
rect 412818 3856 412824 3868
rect 169076 3828 412824 3856
rect 169076 3816 169082 3828
rect 412818 3816 412824 3828
rect 412876 3816 412882 3868
rect 423766 3816 423772 3868
rect 423824 3856 423830 3868
rect 424962 3856 424968 3868
rect 423824 3828 424968 3856
rect 423824 3816 423830 3828
rect 424962 3816 424968 3828
rect 425020 3816 425026 3868
rect 440326 3816 440332 3868
rect 440384 3856 440390 3868
rect 441522 3856 441528 3868
rect 440384 3828 441528 3856
rect 440384 3816 440390 3828
rect 441522 3816 441528 3828
rect 441580 3816 441586 3868
rect 446398 3816 446404 3868
rect 446456 3856 446462 3868
rect 446456 3828 451274 3856
rect 446456 3816 446462 3828
rect 35250 3748 35256 3800
rect 35308 3788 35314 3800
rect 53098 3788 53104 3800
rect 35308 3760 53104 3788
rect 35308 3748 35314 3760
rect 53098 3748 53104 3760
rect 53156 3748 53162 3800
rect 66162 3748 66168 3800
rect 66220 3788 66226 3800
rect 85758 3788 85764 3800
rect 66220 3760 85764 3788
rect 66220 3748 66226 3760
rect 85758 3748 85764 3760
rect 85816 3748 85822 3800
rect 92290 3748 92296 3800
rect 92348 3788 92354 3800
rect 109218 3788 109224 3800
rect 92348 3760 109224 3788
rect 92348 3748 92354 3760
rect 109218 3748 109224 3760
rect 109276 3748 109282 3800
rect 119338 3748 119344 3800
rect 119396 3788 119402 3800
rect 126882 3788 126888 3800
rect 119396 3760 126888 3788
rect 119396 3748 119402 3760
rect 126882 3748 126888 3760
rect 126940 3748 126946 3800
rect 127894 3748 127900 3800
rect 127952 3788 127958 3800
rect 442626 3788 442632 3800
rect 127952 3760 442632 3788
rect 127952 3748 127958 3760
rect 442626 3748 442632 3760
rect 442684 3748 442690 3800
rect 445846 3748 445852 3800
rect 445904 3788 445910 3800
rect 447042 3788 447048 3800
rect 445904 3760 447048 3788
rect 445904 3748 445910 3760
rect 447042 3748 447048 3760
rect 447100 3748 447106 3800
rect 451246 3788 451274 3828
rect 523218 3788 523224 3800
rect 451246 3760 523224 3788
rect 523218 3748 523224 3760
rect 523276 3748 523282 3800
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 83918 3720 83924 3732
rect 41932 3692 83924 3720
rect 41932 3680 41938 3692
rect 83918 3680 83924 3692
rect 83976 3680 83982 3732
rect 88610 3680 88616 3732
rect 88668 3720 88674 3732
rect 102594 3720 102600 3732
rect 88668 3692 102600 3720
rect 88668 3680 88674 3692
rect 102594 3680 102600 3692
rect 102652 3680 102658 3732
rect 104434 3680 104440 3732
rect 104492 3720 104498 3732
rect 123570 3720 123576 3732
rect 104492 3692 123576 3720
rect 104492 3680 104498 3692
rect 123570 3680 123576 3692
rect 123628 3680 123634 3732
rect 128078 3680 128084 3732
rect 128136 3720 128142 3732
rect 456702 3720 456708 3732
rect 128136 3692 456708 3720
rect 128136 3680 128142 3692
rect 456702 3680 456708 3692
rect 456760 3680 456766 3732
rect 456886 3680 456892 3732
rect 456944 3720 456950 3732
rect 458082 3720 458088 3732
rect 456944 3692 458088 3720
rect 456944 3680 456950 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 462406 3680 462412 3732
rect 462464 3720 462470 3732
rect 463602 3720 463608 3732
rect 462464 3692 463608 3720
rect 462464 3680 462470 3692
rect 463602 3680 463608 3692
rect 463660 3680 463666 3732
rect 476850 3720 476856 3732
rect 470566 3692 476856 3720
rect 37458 3612 37464 3664
rect 37516 3652 37522 3664
rect 83090 3652 83096 3664
rect 37516 3624 83096 3652
rect 37516 3612 37522 3624
rect 83090 3612 83096 3624
rect 83148 3612 83154 3664
rect 92106 3612 92112 3664
rect 92164 3652 92170 3664
rect 125778 3652 125784 3664
rect 92164 3624 125784 3652
rect 92164 3612 92170 3624
rect 125778 3612 125784 3624
rect 125836 3612 125842 3664
rect 127986 3612 127992 3664
rect 128044 3652 128050 3664
rect 470566 3652 470594 3692
rect 476850 3680 476856 3692
rect 476908 3680 476914 3732
rect 473538 3652 473544 3664
rect 128044 3624 470594 3652
rect 473372 3624 473544 3652
rect 128044 3612 128050 3624
rect 33042 3544 33048 3596
rect 33100 3584 33106 3596
rect 75730 3584 75736 3596
rect 33100 3556 75736 3584
rect 33100 3544 33106 3556
rect 75730 3544 75736 3556
rect 75788 3544 75794 3596
rect 80054 3584 80060 3596
rect 75840 3556 80060 3584
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 31018 3516 31024 3528
rect 27580 3488 31024 3516
rect 27580 3476 27586 3488
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 75840 3516 75868 3556
rect 80054 3544 80060 3556
rect 80112 3544 80118 3596
rect 87322 3584 87328 3596
rect 84166 3556 87328 3584
rect 32324 3488 75868 3516
rect 29730 3408 29736 3460
rect 29788 3448 29794 3460
rect 32324 3448 32352 3488
rect 75914 3476 75920 3528
rect 75972 3516 75978 3528
rect 77202 3516 77208 3528
rect 75972 3488 77208 3516
rect 75972 3476 75978 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 82722 3476 82728 3528
rect 82780 3516 82786 3528
rect 84166 3516 84194 3556
rect 87322 3544 87328 3556
rect 87380 3544 87386 3596
rect 90726 3544 90732 3596
rect 90784 3584 90790 3596
rect 90784 3556 91692 3584
rect 90784 3544 90790 3556
rect 82780 3488 84194 3516
rect 82780 3476 82786 3488
rect 86034 3476 86040 3528
rect 86092 3516 86098 3528
rect 87230 3516 87236 3528
rect 86092 3488 87236 3516
rect 86092 3476 86098 3488
rect 87230 3476 87236 3488
rect 87288 3476 87294 3528
rect 89346 3476 89352 3528
rect 89404 3516 89410 3528
rect 91554 3516 91560 3528
rect 89404 3488 91560 3516
rect 89404 3476 89410 3488
rect 91554 3476 91560 3488
rect 91612 3476 91618 3528
rect 91664 3516 91692 3556
rect 91922 3544 91928 3596
rect 91980 3584 91986 3596
rect 112530 3584 112536 3596
rect 91980 3556 112536 3584
rect 91980 3544 91986 3556
rect 112530 3544 112536 3556
rect 112588 3544 112594 3596
rect 121270 3544 121276 3596
rect 121328 3584 121334 3596
rect 473372 3584 473400 3624
rect 473538 3612 473544 3624
rect 473596 3612 473602 3664
rect 121328 3556 473400 3584
rect 121328 3544 121334 3556
rect 473446 3544 473452 3596
rect 473504 3584 473510 3596
rect 474642 3584 474648 3596
rect 473504 3556 474648 3584
rect 473504 3544 473510 3556
rect 474642 3544 474648 3556
rect 474700 3544 474706 3596
rect 484394 3544 484400 3596
rect 484452 3584 484458 3596
rect 485682 3584 485688 3596
rect 484452 3556 485688 3584
rect 484452 3544 484458 3556
rect 485682 3544 485688 3556
rect 485740 3544 485746 3596
rect 493410 3584 493416 3596
rect 489886 3556 493416 3584
rect 115842 3516 115848 3528
rect 91664 3488 115848 3516
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 122558 3476 122564 3528
rect 122616 3516 122622 3528
rect 489886 3516 489914 3556
rect 493410 3544 493416 3556
rect 493468 3544 493474 3596
rect 501046 3544 501052 3596
rect 501104 3584 501110 3596
rect 502242 3584 502248 3596
rect 501104 3556 502248 3584
rect 501104 3544 501110 3556
rect 502242 3544 502248 3556
rect 502300 3544 502306 3596
rect 506566 3544 506572 3596
rect 506624 3584 506630 3596
rect 507762 3584 507768 3596
rect 506624 3556 507768 3584
rect 506624 3544 506630 3556
rect 507762 3544 507768 3556
rect 507820 3544 507826 3596
rect 545206 3544 545212 3596
rect 545264 3584 545270 3596
rect 546402 3584 546408 3596
rect 545264 3556 546408 3584
rect 545264 3544 545270 3556
rect 546402 3544 546408 3556
rect 546460 3544 546466 3596
rect 550726 3544 550732 3596
rect 550784 3584 550790 3596
rect 551922 3584 551928 3596
rect 550784 3556 551928 3584
rect 550784 3544 550790 3556
rect 551922 3544 551928 3556
rect 551980 3544 551986 3596
rect 122616 3488 489914 3516
rect 122616 3476 122622 3488
rect 490006 3476 490012 3528
rect 490064 3516 490070 3528
rect 491202 3516 491208 3528
rect 490064 3488 491208 3516
rect 490064 3476 490070 3488
rect 491202 3476 491208 3488
rect 491260 3476 491266 3528
rect 511994 3476 512000 3528
rect 512052 3516 512058 3528
rect 513282 3516 513288 3528
rect 512052 3488 513288 3516
rect 512052 3476 512058 3488
rect 513282 3476 513288 3488
rect 513340 3476 513346 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540882 3516 540888 3528
rect 539652 3488 540888 3516
rect 539652 3476 539658 3488
rect 540882 3476 540888 3488
rect 540940 3476 540946 3528
rect 82998 3448 83004 3460
rect 29788 3420 32352 3448
rect 35866 3420 83004 3448
rect 29788 3408 29794 3420
rect 28626 3340 28632 3392
rect 28684 3380 28690 3392
rect 35866 3380 35894 3420
rect 82998 3408 83004 3420
rect 83056 3408 83062 3460
rect 87414 3408 87420 3460
rect 87472 3448 87478 3460
rect 90450 3448 90456 3460
rect 87472 3420 90456 3448
rect 87472 3408 87478 3420
rect 90450 3408 90456 3420
rect 90508 3408 90514 3460
rect 118050 3448 118056 3460
rect 93826 3420 118056 3448
rect 28684 3352 35894 3380
rect 28684 3340 28690 3352
rect 59354 3340 59360 3392
rect 59412 3380 59418 3392
rect 60642 3380 60648 3392
rect 59412 3352 60648 3380
rect 59412 3340 59418 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 70394 3340 70400 3392
rect 70452 3380 70458 3392
rect 71682 3380 71688 3392
rect 70452 3352 71688 3380
rect 70452 3340 70458 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 88518 3340 88524 3392
rect 88576 3380 88582 3392
rect 92658 3380 92664 3392
rect 88576 3352 92664 3380
rect 88576 3340 88582 3352
rect 92658 3340 92664 3352
rect 92716 3340 92722 3392
rect 89806 3272 89812 3324
rect 89864 3312 89870 3324
rect 93826 3312 93854 3420
rect 118050 3408 118056 3420
rect 118108 3408 118114 3460
rect 121546 3408 121552 3460
rect 121604 3448 121610 3460
rect 496722 3448 496728 3460
rect 121604 3420 496728 3448
rect 121604 3408 121610 3420
rect 496722 3408 496728 3420
rect 496780 3408 496786 3460
rect 100018 3340 100024 3392
rect 100076 3380 100082 3392
rect 101490 3380 101496 3392
rect 100076 3352 101496 3380
rect 100076 3340 100082 3352
rect 101490 3340 101496 3352
rect 101548 3340 101554 3392
rect 135898 3340 135904 3392
rect 135956 3380 135962 3392
rect 137922 3380 137928 3392
rect 135956 3352 137928 3380
rect 135956 3340 135962 3352
rect 137922 3340 137928 3352
rect 137980 3340 137986 3392
rect 153194 3340 153200 3392
rect 153252 3380 153258 3392
rect 154482 3380 154488 3392
rect 153252 3352 154488 3380
rect 153252 3340 153258 3352
rect 154482 3340 154488 3352
rect 154540 3340 154546 3392
rect 164142 3340 164148 3392
rect 164200 3380 164206 3392
rect 167730 3380 167736 3392
rect 164200 3352 167736 3380
rect 164200 3340 164206 3352
rect 167730 3340 167736 3352
rect 167788 3340 167794 3392
rect 180794 3340 180800 3392
rect 180852 3380 180858 3392
rect 182082 3380 182088 3392
rect 180852 3352 182088 3380
rect 180852 3340 180858 3352
rect 182082 3340 182088 3352
rect 182140 3340 182146 3392
rect 186314 3340 186320 3392
rect 186372 3380 186378 3392
rect 187602 3380 187608 3392
rect 186372 3352 187608 3380
rect 186372 3340 186378 3352
rect 187602 3340 187608 3352
rect 187660 3340 187666 3392
rect 197354 3340 197360 3392
rect 197412 3380 197418 3392
rect 198642 3380 198648 3392
rect 197412 3352 198648 3380
rect 197412 3340 197418 3352
rect 198642 3340 198648 3352
rect 198700 3340 198706 3392
rect 202874 3340 202880 3392
rect 202932 3380 202938 3392
rect 204162 3380 204168 3392
rect 202932 3352 204168 3380
rect 202932 3340 202938 3352
rect 204162 3340 204168 3352
rect 204220 3340 204226 3392
rect 235994 3340 236000 3392
rect 236052 3380 236058 3392
rect 237282 3380 237288 3392
rect 236052 3352 237288 3380
rect 236052 3340 236058 3352
rect 237282 3340 237288 3352
rect 237340 3340 237346 3392
rect 252554 3340 252560 3392
rect 252612 3380 252618 3392
rect 253842 3380 253848 3392
rect 252612 3352 253848 3380
rect 252612 3340 252618 3352
rect 253842 3340 253848 3352
rect 253900 3340 253906 3392
rect 269114 3340 269120 3392
rect 269172 3380 269178 3392
rect 270402 3380 270408 3392
rect 269172 3352 270408 3380
rect 269172 3340 269178 3352
rect 270402 3340 270408 3352
rect 270460 3340 270466 3392
rect 285674 3340 285680 3392
rect 285732 3380 285738 3392
rect 286962 3380 286968 3392
rect 285732 3352 286968 3380
rect 285732 3340 285738 3352
rect 286962 3340 286968 3352
rect 287020 3340 287026 3392
rect 302234 3340 302240 3392
rect 302292 3380 302298 3392
rect 303522 3380 303528 3392
rect 302292 3352 303528 3380
rect 302292 3340 302298 3352
rect 303522 3340 303528 3352
rect 303580 3340 303586 3392
rect 313274 3340 313280 3392
rect 313332 3380 313338 3392
rect 314562 3380 314568 3392
rect 313332 3352 314568 3380
rect 313332 3340 313338 3352
rect 314562 3340 314568 3352
rect 314620 3340 314626 3392
rect 318794 3340 318800 3392
rect 318852 3380 318858 3392
rect 320082 3380 320088 3392
rect 318852 3352 320088 3380
rect 318852 3340 318858 3352
rect 320082 3340 320088 3352
rect 320140 3340 320146 3392
rect 335354 3340 335360 3392
rect 335412 3380 335418 3392
rect 336642 3380 336648 3392
rect 335412 3352 336648 3380
rect 335412 3340 335418 3352
rect 336642 3340 336648 3352
rect 336700 3340 336706 3392
rect 351914 3340 351920 3392
rect 351972 3380 351978 3392
rect 353202 3380 353208 3392
rect 351972 3352 353208 3380
rect 351972 3340 351978 3352
rect 353202 3340 353208 3352
rect 353260 3340 353266 3392
rect 362954 3340 362960 3392
rect 363012 3380 363018 3392
rect 364242 3380 364248 3392
rect 363012 3352 364248 3380
rect 363012 3340 363018 3352
rect 364242 3340 364248 3352
rect 364300 3340 364306 3392
rect 368474 3340 368480 3392
rect 368532 3380 368538 3392
rect 369762 3380 369768 3392
rect 368532 3352 369768 3380
rect 368532 3340 368538 3352
rect 369762 3340 369768 3352
rect 369820 3340 369826 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 379514 3340 379520 3392
rect 379572 3380 379578 3392
rect 380802 3380 380808 3392
rect 379572 3352 380808 3380
rect 379572 3340 379578 3352
rect 380802 3340 380808 3352
rect 380860 3340 380866 3392
rect 385034 3340 385040 3392
rect 385092 3380 385098 3392
rect 386322 3380 386328 3392
rect 385092 3352 386328 3380
rect 385092 3340 385098 3352
rect 386322 3340 386328 3352
rect 386380 3340 386386 3392
rect 401594 3340 401600 3392
rect 401652 3380 401658 3392
rect 402882 3380 402888 3392
rect 401652 3352 402888 3380
rect 401652 3340 401658 3352
rect 402882 3340 402888 3352
rect 402940 3340 402946 3392
rect 412726 3340 412732 3392
rect 412784 3380 412790 3392
rect 413922 3380 413928 3392
rect 412784 3352 413928 3380
rect 412784 3340 412790 3352
rect 413922 3340 413928 3352
rect 413980 3340 413986 3392
rect 418154 3340 418160 3392
rect 418212 3380 418218 3392
rect 419442 3380 419448 3392
rect 418212 3352 419448 3380
rect 418212 3340 418218 3352
rect 419442 3340 419448 3352
rect 419500 3340 419506 3392
rect 429194 3340 429200 3392
rect 429252 3380 429258 3392
rect 430482 3380 430488 3392
rect 429252 3352 430488 3380
rect 429252 3340 429258 3352
rect 430482 3340 430488 3352
rect 430540 3340 430546 3392
rect 434714 3340 434720 3392
rect 434772 3380 434778 3392
rect 436002 3380 436008 3392
rect 434772 3352 436008 3380
rect 434772 3340 434778 3352
rect 436002 3340 436008 3352
rect 436060 3340 436066 3392
rect 451274 3340 451280 3392
rect 451332 3380 451338 3392
rect 452562 3380 452568 3392
rect 451332 3352 452568 3380
rect 451332 3340 451338 3352
rect 452562 3340 452568 3352
rect 452620 3340 452626 3392
rect 456702 3340 456708 3392
rect 456760 3380 456766 3392
rect 459186 3380 459192 3392
rect 456760 3352 459192 3380
rect 456760 3340 456766 3352
rect 459186 3340 459192 3352
rect 459244 3340 459250 3392
rect 89864 3284 93854 3312
rect 89864 3272 89870 3284
rect 131758 3204 131764 3256
rect 131816 3244 131822 3256
rect 133506 3244 133512 3256
rect 131816 3216 133512 3244
rect 131816 3204 131822 3216
rect 133506 3204 133512 3216
rect 133564 3204 133570 3256
rect 87138 3136 87144 3188
rect 87196 3176 87202 3188
rect 89346 3176 89352 3188
rect 87196 3148 89352 3176
rect 87196 3136 87202 3148
rect 89346 3136 89352 3148
rect 89404 3136 89410 3188
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 43438 3040 43444 3052
rect 36412 3012 43444 3040
rect 36412 3000 36418 3012
rect 43438 3000 43444 3012
rect 43496 3000 43502 3052
rect 80514 2796 80520 2848
rect 80572 2836 80578 2848
rect 82354 2836 82360 2848
rect 80572 2808 82360 2836
rect 80572 2796 80578 2808
rect 82354 2796 82360 2808
rect 82412 2796 82418 2848
rect 478874 1096 478880 1148
rect 478932 1136 478938 1148
rect 480162 1136 480168 1148
rect 478932 1108 480168 1136
rect 478932 1096 478938 1108
rect 480162 1096 480168 1108
rect 480220 1096 480226 1148
rect 534074 688 534080 740
rect 534132 728 534138 740
rect 535362 728 535368 740
rect 534132 700 535368 728
rect 534132 688 534138 700
rect 535362 688 535368 700
rect 535420 688 535426 740
<< via1 >>
rect 74540 702992 74592 703044
rect 75736 702992 75788 703044
rect 204260 702992 204312 703044
rect 205456 702992 205508 703044
rect 333980 702992 334032 703044
rect 335176 702992 335228 703044
rect 463700 702992 463752 703044
rect 464896 702992 464948 703044
rect 97356 700748 97408 700800
rect 109040 700748 109092 700800
rect 107660 700680 107712 700732
rect 162216 700680 162268 700732
rect 32496 700612 32548 700664
rect 110972 700612 111024 700664
rect 107752 700544 107804 700596
rect 227076 700544 227128 700596
rect 106280 700476 106332 700528
rect 291936 700476 291988 700528
rect 103520 700408 103572 700460
rect 421656 700408 421708 700460
rect 102140 700340 102192 700392
rect 486516 700340 486568 700392
rect 102232 700272 102284 700324
rect 551376 700272 551428 700324
rect 100852 695512 100904 695564
rect 580172 695512 580224 695564
rect 3424 694152 3476 694204
rect 111248 694152 111300 694204
rect 101036 680348 101088 680400
rect 580172 680348 580224 680400
rect 3424 677560 3476 677612
rect 112168 677560 112220 677612
rect 100208 663756 100260 663808
rect 580172 663756 580224 663808
rect 3424 661036 3476 661088
rect 111892 661036 111944 661088
rect 99656 648592 99708 648644
rect 580172 648592 580224 648644
rect 3240 644444 3292 644496
rect 112352 644444 112404 644496
rect 99932 633428 99984 633480
rect 580172 633428 580224 633480
rect 3424 627920 3476 627972
rect 113364 627920 113416 627972
rect 99472 616836 99524 616888
rect 580172 616836 580224 616888
rect 3424 609968 3476 610020
rect 111064 609968 111116 610020
rect 98552 601672 98604 601724
rect 580172 601672 580224 601724
rect 98276 586508 98328 586560
rect 580908 586508 580960 586560
rect 3056 576852 3108 576904
rect 114008 576852 114060 576904
rect 98368 569916 98420 569968
rect 580172 569916 580224 569968
rect 3056 560260 3108 560312
rect 112444 560260 112496 560312
rect 97448 554752 97500 554804
rect 580172 554752 580224 554804
rect 96896 539588 96948 539640
rect 580172 539588 580224 539640
rect 3608 527144 3660 527196
rect 115112 527144 115164 527196
rect 97172 522996 97224 523048
rect 580172 522996 580224 523048
rect 3332 510620 3384 510672
rect 112536 510620 112588 510672
rect 95792 507832 95844 507884
rect 580172 507832 580224 507884
rect 3332 494028 3384 494080
rect 116492 494028 116544 494080
rect 96712 492668 96764 492720
rect 580172 492668 580224 492720
rect 3148 476144 3200 476196
rect 116768 476144 116820 476196
rect 95516 476076 95568 476128
rect 580172 476076 580224 476128
rect 95332 460912 95384 460964
rect 580172 460912 580224 460964
rect 3148 459552 3200 459604
rect 113824 459552 113876 459604
rect 95608 445748 95660 445800
rect 580172 445748 580224 445800
rect 3332 442960 3384 443012
rect 117044 442960 117096 443012
rect 94688 429156 94740 429208
rect 580172 429156 580224 429208
rect 3332 426436 3384 426488
rect 117596 426436 117648 426488
rect 94136 413992 94188 414044
rect 580172 413992 580224 414044
rect 3332 409844 3384 409896
rect 113916 409844 113968 409896
rect 94412 398828 94464 398880
rect 580172 398828 580224 398880
rect 3608 393320 3660 393372
rect 117872 393320 117924 393372
rect 93952 382236 94004 382288
rect 580172 382236 580224 382288
rect 3332 376728 3384 376780
rect 117964 376728 118016 376780
rect 92480 367072 92532 367124
rect 580172 367072 580224 367124
rect 3332 360204 3384 360256
rect 115204 360204 115256 360256
rect 92756 351908 92808 351960
rect 580172 351908 580224 351960
rect 3332 342252 3384 342304
rect 119344 342252 119396 342304
rect 92848 335316 92900 335368
rect 580172 335316 580224 335368
rect 3332 325660 3384 325712
rect 118056 325660 118108 325712
rect 91100 320152 91152 320204
rect 580172 320152 580224 320204
rect 3332 309136 3384 309188
rect 119620 309136 119672 309188
rect 91376 304988 91428 305040
rect 580172 304988 580224 305040
rect 3332 292544 3384 292596
rect 120632 292544 120684 292596
rect 91652 288396 91704 288448
rect 580172 288396 580224 288448
rect 3332 276020 3384 276072
rect 120724 276020 120776 276072
rect 89720 273232 89772 273284
rect 580172 273232 580224 273284
rect 2964 259428 3016 259480
rect 120448 259428 120500 259480
rect 91192 258068 91244 258120
rect 580908 258068 580960 258120
rect 3332 242904 3384 242956
rect 120356 242904 120408 242956
rect 89996 241476 90048 241528
rect 580172 241476 580224 241528
rect 3332 226380 3384 226432
rect 118148 226380 118200 226432
rect 89812 226312 89864 226364
rect 580172 226312 580224 226364
rect 90088 211148 90140 211200
rect 580172 211148 580224 211200
rect 3332 209788 3384 209840
rect 116584 209788 116636 209840
rect 88340 194556 88392 194608
rect 580172 194556 580224 194608
rect 3332 191836 3384 191888
rect 121736 191836 121788 191888
rect 88616 179392 88668 179444
rect 580172 179392 580224 179444
rect 3056 175244 3108 175296
rect 122012 175244 122064 175296
rect 88892 164228 88944 164280
rect 580172 164228 580224 164280
rect 88340 160216 88392 160268
rect 89444 160216 89496 160268
rect 92756 159196 92808 159248
rect 93308 159196 93360 159248
rect 107660 158856 107712 158908
rect 108764 158856 108816 158908
rect 3148 158720 3200 158772
rect 116492 158720 116544 158772
rect 102140 158244 102192 158296
rect 103244 158244 103296 158296
rect 108488 157020 108540 157072
rect 139400 157020 139452 157072
rect 74540 156952 74592 157004
rect 109684 156952 109736 157004
rect 107384 156884 107436 156936
rect 204260 156884 204312 156936
rect 9680 156816 9732 156868
rect 110696 156816 110748 156868
rect 120356 156816 120408 156868
rect 120908 156816 120960 156868
rect 106372 156748 106424 156800
rect 269120 156748 269172 156800
rect 105084 156680 105136 156732
rect 333980 156680 334032 156732
rect 105452 156612 105504 156664
rect 356060 156612 356112 156664
rect 120356 156544 120408 156596
rect 120632 156544 120684 156596
rect 113916 155864 113968 155916
rect 117504 155864 117556 155916
rect 118056 155864 118108 155916
rect 119804 155864 119856 155916
rect 108212 155592 108264 155644
rect 183560 155592 183612 155644
rect 3424 155524 3476 155576
rect 113732 155524 113784 155576
rect 3516 155456 3568 155508
rect 114928 155456 114980 155508
rect 107108 155388 107160 155440
rect 248420 155388 248472 155440
rect 104072 155320 104124 155372
rect 398840 155320 398892 155372
rect 102968 155252 103020 155304
rect 463700 155252 463752 155304
rect 101864 155184 101916 155236
rect 528560 155184 528612 155236
rect 117964 154504 118016 154556
rect 118700 154504 118752 154556
rect 109592 154232 109644 154284
rect 118792 154232 118844 154284
rect 53840 154164 53892 154216
rect 110420 154164 110472 154216
rect 106188 154096 106240 154148
rect 313280 154096 313332 154148
rect 104992 154028 105044 154080
rect 378140 154028 378192 154080
rect 103980 153960 104032 154012
rect 443000 153960 443052 154012
rect 102876 153892 102928 153944
rect 507860 153892 507912 153944
rect 101772 153824 101824 153876
rect 572720 153824 572772 153876
rect 89996 153280 90048 153332
rect 90548 153280 90600 153332
rect 91376 153280 91428 153332
rect 92204 153280 92256 153332
rect 92480 153280 92532 153332
rect 93032 153280 93084 153332
rect 95516 153280 95568 153332
rect 96068 153280 96120 153332
rect 96896 153280 96948 153332
rect 97724 153280 97776 153332
rect 98276 153280 98328 153332
rect 98828 153280 98880 153332
rect 89720 153212 89772 153264
rect 90824 153212 90876 153264
rect 91100 153212 91152 153264
rect 91928 153212 91980 153264
rect 111064 153144 111116 153196
rect 112904 153144 112956 153196
rect 113824 153144 113876 153196
rect 116308 153144 116360 153196
rect 118148 153144 118200 153196
rect 121460 153144 121512 153196
rect 115204 153076 115256 153128
rect 118424 153076 118476 153128
rect 116584 153008 116636 153060
rect 121184 153008 121236 153060
rect 116492 152940 116544 152992
rect 122012 152940 122064 152992
rect 109316 152872 109368 152924
rect 128728 152872 128780 152924
rect 7564 152668 7616 152720
rect 123116 152804 123168 152856
rect 81900 152532 81952 152584
rect 95792 152532 95844 152584
rect 80888 152464 80940 152516
rect 94688 152464 94740 152516
rect 114836 152464 114888 152516
rect 118056 152464 118108 152516
rect 4804 152396 4856 152448
rect 122840 152668 122892 152720
rect 3792 152328 3844 152380
rect 123944 152328 123996 152380
rect 82360 152260 82412 152312
rect 101312 152260 101364 152312
rect 115848 152260 115900 152312
rect 127992 152260 128044 152312
rect 82176 152192 82228 152244
rect 96896 152192 96948 152244
rect 108120 152192 108172 152244
rect 81716 152124 81768 152176
rect 99104 152124 99156 152176
rect 111432 152124 111484 152176
rect 117780 152124 117832 152176
rect 118056 152192 118108 152244
rect 128544 152192 128596 152244
rect 128452 152124 128504 152176
rect 81440 152056 81492 152108
rect 100208 152056 100260 152108
rect 104808 152056 104860 152108
rect 128360 152056 128412 152108
rect 85856 151988 85908 152040
rect 95240 151988 95292 152040
rect 103796 151988 103848 152040
rect 128820 151988 128872 152040
rect 113640 151920 113692 151972
rect 128912 151920 128964 151972
rect 112444 151852 112496 151904
rect 114008 151852 114060 151904
rect 117780 151852 117832 151904
rect 128636 151852 128688 151904
rect 82268 151784 82320 151836
rect 98184 151784 98236 151836
rect 112536 151784 112588 151836
rect 115020 151784 115072 151836
rect 116952 151784 117004 151836
rect 128176 151784 128228 151836
rect 3516 151104 3568 151156
rect 98000 151104 98052 151156
rect 95240 151036 95292 151088
rect 580356 151036 580408 151088
rect 87788 150764 87840 150816
rect 129004 150764 129056 150816
rect 3884 150696 3936 150748
rect 123392 150696 123444 150748
rect 3700 150628 3752 150680
rect 123668 150628 123720 150680
rect 3608 150560 3660 150612
rect 124220 150560 124272 150612
rect 3240 150492 3292 150544
rect 124496 150492 124548 150544
rect 88524 150424 88576 150476
rect 580172 150424 580224 150476
rect 80980 150152 81032 150204
rect 91514 150152 91566 150204
rect 81348 149948 81400 150000
rect 81164 149880 81216 149932
rect 81072 149744 81124 149796
rect 93584 149812 93636 149864
rect 112352 149812 112404 149864
rect 112628 149812 112680 149864
rect 81256 149676 81308 149728
rect 89168 149676 89220 149728
rect 90272 149744 90324 149796
rect 92480 149676 92532 149728
rect 85304 149608 85356 149660
rect 89444 149608 89496 149660
rect 91652 149608 91704 149660
rect 81808 149540 81860 149592
rect 86960 149540 87012 149592
rect 91928 149540 91980 149592
rect 81992 149472 82044 149524
rect 85856 149472 85908 149524
rect 82084 149404 82136 149456
rect 84568 149404 84620 149456
rect 3424 149336 3476 149388
rect 86408 149404 86460 149456
rect 86684 149472 86736 149524
rect 89444 149404 89496 149456
rect 91652 149404 91704 149456
rect 91928 149404 91980 149456
rect 94136 149404 94188 149456
rect 118148 149540 118200 149592
rect 128084 149540 128136 149592
rect 122564 149404 122616 149456
rect 580264 149404 580316 149456
rect 580632 149268 580684 149320
rect 580540 149200 580592 149252
rect 580448 149132 580500 149184
rect 129004 133832 129056 133884
rect 579988 133832 580040 133884
rect 3332 126420 3384 126472
rect 7564 126420 7616 126472
rect 138664 118600 138716 118652
rect 580172 118600 580224 118652
rect 2780 110100 2832 110152
rect 4804 110100 4856 110152
rect 81900 101464 81952 101516
rect 82360 101464 82412 101516
rect 81808 100240 81860 100292
rect 80888 100172 80940 100224
rect 81808 100104 81860 100156
rect 77852 100036 77904 100088
rect 80428 99968 80480 100020
rect 86638 100104 86690 100156
rect 81440 99900 81492 99952
rect 82360 99900 82412 99952
rect 81624 99832 81676 99884
rect 82590 99832 82642 99884
rect 81440 99764 81492 99816
rect 81900 99764 81952 99816
rect 79784 99696 79836 99748
rect 83510 99900 83562 99952
rect 83602 99900 83654 99952
rect 84062 99900 84114 99952
rect 84154 99900 84206 99952
rect 84246 99900 84298 99952
rect 84338 99900 84390 99952
rect 82774 99832 82826 99884
rect 83050 99832 83102 99884
rect 83326 99832 83378 99884
rect 82912 99628 82964 99680
rect 83234 99764 83286 99816
rect 83188 99628 83240 99680
rect 83786 99764 83838 99816
rect 83556 99628 83608 99680
rect 83648 99628 83700 99680
rect 83372 99492 83424 99544
rect 83832 99492 83884 99544
rect 84614 99832 84666 99884
rect 84706 99832 84758 99884
rect 84384 99764 84436 99816
rect 84200 99696 84252 99748
rect 84476 99628 84528 99680
rect 84476 99492 84528 99544
rect 84568 99424 84620 99476
rect 84660 99424 84712 99476
rect 85166 99900 85218 99952
rect 85994 99900 86046 99952
rect 86178 99900 86230 99952
rect 86270 99900 86322 99952
rect 85810 99832 85862 99884
rect 85902 99832 85954 99884
rect 85350 99764 85402 99816
rect 85626 99764 85678 99816
rect 85396 99628 85448 99680
rect 85672 99628 85724 99680
rect 85304 99560 85356 99612
rect 86040 99628 86092 99680
rect 84936 99424 84988 99476
rect 85212 99424 85264 99476
rect 86592 99832 86644 99884
rect 86316 99764 86368 99816
rect 86454 99764 86506 99816
rect 86730 99764 86782 99816
rect 86592 99696 86644 99748
rect 86776 99628 86828 99680
rect 86408 99560 86460 99612
rect 86684 99424 86736 99476
rect 87006 99900 87058 99952
rect 87834 99900 87886 99952
rect 88018 99900 88070 99952
rect 88478 99900 88530 99952
rect 88570 99900 88622 99952
rect 87558 99832 87610 99884
rect 87190 99764 87242 99816
rect 87282 99764 87334 99816
rect 87144 99560 87196 99612
rect 87512 99696 87564 99748
rect 87880 99628 87932 99680
rect 87788 99560 87840 99612
rect 87420 99492 87472 99544
rect 87604 99492 87656 99544
rect 84844 99356 84896 99408
rect 86224 99356 86276 99408
rect 87052 99288 87104 99340
rect 87880 99492 87932 99544
rect 88294 99832 88346 99884
rect 88340 99628 88392 99680
rect 88156 99560 88208 99612
rect 88432 99424 88484 99476
rect 88754 99832 88806 99884
rect 88938 99900 88990 99952
rect 89214 99900 89266 99952
rect 89306 99900 89358 99952
rect 89582 99900 89634 99952
rect 89168 99696 89220 99748
rect 88984 99628 89036 99680
rect 89490 99764 89542 99816
rect 89444 99628 89496 99680
rect 89536 99628 89588 99680
rect 89076 99492 89128 99544
rect 89904 99492 89956 99544
rect 88708 99424 88760 99476
rect 89352 99356 89404 99408
rect 90502 100036 90554 100088
rect 93722 100036 93774 100088
rect 90318 99900 90370 99952
rect 90410 99900 90462 99952
rect 90594 99900 90646 99952
rect 90226 99832 90278 99884
rect 90364 99696 90416 99748
rect 90640 99764 90692 99816
rect 90548 99628 90600 99680
rect 91238 99900 91290 99952
rect 91330 99764 91382 99816
rect 91008 99560 91060 99612
rect 91192 99628 91244 99680
rect 91284 99560 91336 99612
rect 90732 99424 90784 99476
rect 90824 99356 90876 99408
rect 91790 99900 91842 99952
rect 92342 99900 92394 99952
rect 92710 99900 92762 99952
rect 92894 99900 92946 99952
rect 92986 99900 93038 99952
rect 93262 99900 93314 99952
rect 93354 99900 93406 99952
rect 91514 99832 91566 99884
rect 91606 99832 91658 99884
rect 92158 99832 92210 99884
rect 91652 99560 91704 99612
rect 92020 99560 92072 99612
rect 92434 99832 92486 99884
rect 92296 99628 92348 99680
rect 92848 99696 92900 99748
rect 93308 99764 93360 99816
rect 93400 99628 93452 99680
rect 93906 99900 93958 99952
rect 93998 99900 94050 99952
rect 93860 99628 93912 99680
rect 92480 99560 92532 99612
rect 93124 99560 93176 99612
rect 93216 99560 93268 99612
rect 93952 99560 94004 99612
rect 97586 100172 97638 100224
rect 94366 99900 94418 99952
rect 94642 99900 94694 99952
rect 94734 99900 94786 99952
rect 94918 99900 94970 99952
rect 95746 99900 95798 99952
rect 95930 99900 95982 99952
rect 96022 99900 96074 99952
rect 96298 99900 96350 99952
rect 96574 99900 96626 99952
rect 92296 99492 92348 99544
rect 94044 99492 94096 99544
rect 94228 99492 94280 99544
rect 94550 99832 94602 99884
rect 94688 99764 94740 99816
rect 95102 99832 95154 99884
rect 94872 99696 94924 99748
rect 95194 99764 95246 99816
rect 94964 99628 95016 99680
rect 93308 99424 93360 99476
rect 93584 99424 93636 99476
rect 95056 99424 95108 99476
rect 95148 99424 95200 99476
rect 93584 99288 93636 99340
rect 81716 99220 81768 99272
rect 95976 99764 96028 99816
rect 95884 99628 95936 99680
rect 96942 99900 96994 99952
rect 96850 99832 96902 99884
rect 96712 99628 96764 99680
rect 97126 99832 97178 99884
rect 97310 99832 97362 99884
rect 96896 99696 96948 99748
rect 97080 99696 97132 99748
rect 97172 99628 97224 99680
rect 97678 99900 97730 99952
rect 97770 99832 97822 99884
rect 97632 99628 97684 99680
rect 97448 99560 97500 99612
rect 97540 99560 97592 99612
rect 97954 99900 98006 99952
rect 98230 99900 98282 99952
rect 98414 99900 98466 99952
rect 98138 99764 98190 99816
rect 98000 99560 98052 99612
rect 96436 99492 96488 99544
rect 97908 99492 97960 99544
rect 98368 99696 98420 99748
rect 98460 99628 98512 99680
rect 98966 100104 99018 100156
rect 128176 100308 128228 100360
rect 99610 100036 99662 100088
rect 98690 99900 98742 99952
rect 98874 99900 98926 99952
rect 99150 99900 99202 99952
rect 99518 99900 99570 99952
rect 99012 99832 99064 99884
rect 99242 99832 99294 99884
rect 99426 99832 99478 99884
rect 99104 99764 99156 99816
rect 98736 99696 98788 99748
rect 98920 99696 98972 99748
rect 98828 99560 98880 99612
rect 99656 99764 99708 99816
rect 99564 99696 99616 99748
rect 99012 99424 99064 99476
rect 100162 99900 100214 99952
rect 100254 99900 100306 99952
rect 100070 99832 100122 99884
rect 99932 99560 99984 99612
rect 99748 99492 99800 99544
rect 100208 99560 100260 99612
rect 99840 99424 99892 99476
rect 100024 99424 100076 99476
rect 100714 100036 100766 100088
rect 104854 100036 104906 100088
rect 107338 100036 107390 100088
rect 112582 100036 112634 100088
rect 100438 99900 100490 99952
rect 100622 99900 100674 99952
rect 100898 99900 100950 99952
rect 101082 99900 101134 99952
rect 101266 99900 101318 99952
rect 101450 99900 101502 99952
rect 101726 99900 101778 99952
rect 100668 99764 100720 99816
rect 100944 99628 100996 99680
rect 101128 99628 101180 99680
rect 101542 99764 101594 99816
rect 101588 99628 101640 99680
rect 100484 99560 100536 99612
rect 101312 99560 101364 99612
rect 101404 99560 101456 99612
rect 101496 99560 101548 99612
rect 100760 99492 100812 99544
rect 101864 99560 101916 99612
rect 102094 99900 102146 99952
rect 102186 99900 102238 99952
rect 102278 99900 102330 99952
rect 102370 99900 102422 99952
rect 102462 99900 102514 99952
rect 102830 99900 102882 99952
rect 102048 99764 102100 99816
rect 101956 99492 102008 99544
rect 101036 99356 101088 99408
rect 102324 99764 102376 99816
rect 102416 99696 102468 99748
rect 102646 99832 102698 99884
rect 103014 99764 103066 99816
rect 102968 99628 103020 99680
rect 102600 99560 102652 99612
rect 102692 99492 102744 99544
rect 103290 99900 103342 99952
rect 103474 99900 103526 99952
rect 103750 99900 103802 99952
rect 103842 99900 103894 99952
rect 103934 99900 103986 99952
rect 104026 99900 104078 99952
rect 104118 99900 104170 99952
rect 103290 99764 103342 99816
rect 103382 99764 103434 99816
rect 103336 99628 103388 99680
rect 103658 99832 103710 99884
rect 103428 99560 103480 99612
rect 103888 99696 103940 99748
rect 103980 99628 104032 99680
rect 104072 99628 104124 99680
rect 103336 99492 103388 99544
rect 103612 99492 103664 99544
rect 103704 99492 103756 99544
rect 103796 99424 103848 99476
rect 104394 99900 104446 99952
rect 104670 99900 104722 99952
rect 104486 99832 104538 99884
rect 104624 99764 104676 99816
rect 104808 99832 104860 99884
rect 105130 99900 105182 99952
rect 105314 99900 105366 99952
rect 105498 99900 105550 99952
rect 106234 99900 106286 99952
rect 106326 99900 106378 99952
rect 106510 99900 106562 99952
rect 106694 99900 106746 99952
rect 105038 99832 105090 99884
rect 104716 99696 104768 99748
rect 104900 99696 104952 99748
rect 104440 99628 104492 99680
rect 104808 99628 104860 99680
rect 105084 99560 105136 99612
rect 102876 99356 102928 99408
rect 104256 99356 104308 99408
rect 105406 99832 105458 99884
rect 105958 99832 106010 99884
rect 106142 99832 106194 99884
rect 106004 99696 106056 99748
rect 106418 99764 106470 99816
rect 106280 99696 106332 99748
rect 105544 99628 105596 99680
rect 106096 99628 106148 99680
rect 106188 99628 106240 99680
rect 106372 99560 106424 99612
rect 105452 99492 105504 99544
rect 106648 99560 106700 99612
rect 106878 99900 106930 99952
rect 106970 99900 107022 99952
rect 107062 99900 107114 99952
rect 106924 99764 106976 99816
rect 107614 99900 107666 99952
rect 107706 99900 107758 99952
rect 107982 99900 108034 99952
rect 108350 99900 108402 99952
rect 108534 99900 108586 99952
rect 109086 99900 109138 99952
rect 107660 99764 107712 99816
rect 107016 99696 107068 99748
rect 107476 99696 107528 99748
rect 107384 99560 107436 99612
rect 108120 99560 108172 99612
rect 106740 99492 106792 99544
rect 108396 99492 108448 99544
rect 108994 99764 109046 99816
rect 108810 99696 108862 99748
rect 109362 99832 109414 99884
rect 109040 99628 109092 99680
rect 108948 99560 109000 99612
rect 108672 99492 108724 99544
rect 106464 99424 106516 99476
rect 108488 99424 108540 99476
rect 109914 99968 109966 100020
rect 109822 99900 109874 99952
rect 110006 99900 110058 99952
rect 110098 99900 110150 99952
rect 110466 99900 110518 99952
rect 109868 99628 109920 99680
rect 110282 99832 110334 99884
rect 110374 99832 110426 99884
rect 110052 99696 110104 99748
rect 110144 99696 110196 99748
rect 110558 99764 110610 99816
rect 110420 99696 110472 99748
rect 110236 99628 110288 99680
rect 110512 99628 110564 99680
rect 110834 99900 110886 99952
rect 111018 99900 111070 99952
rect 111110 99900 111162 99952
rect 111570 99900 111622 99952
rect 111478 99832 111530 99884
rect 111662 99832 111714 99884
rect 111156 99764 111208 99816
rect 111432 99696 111484 99748
rect 111064 99560 111116 99612
rect 109960 99492 110012 99544
rect 110696 99492 110748 99544
rect 110880 99492 110932 99544
rect 111616 99628 111668 99680
rect 112030 99900 112082 99952
rect 111846 99832 111898 99884
rect 111340 99560 111392 99612
rect 111524 99560 111576 99612
rect 111708 99560 111760 99612
rect 109684 99424 109736 99476
rect 106004 99356 106056 99408
rect 96068 99220 96120 99272
rect 111616 99220 111668 99272
rect 111984 99628 112036 99680
rect 111984 99356 112036 99408
rect 112306 99832 112358 99884
rect 117642 100104 117694 100156
rect 113870 99968 113922 100020
rect 113134 99832 113186 99884
rect 113272 99628 113324 99680
rect 113686 99900 113738 99952
rect 114146 99900 114198 99952
rect 113502 99832 113554 99884
rect 113640 99628 113692 99680
rect 113824 99628 113876 99680
rect 113916 99628 113968 99680
rect 114100 99628 114152 99680
rect 113456 99560 113508 99612
rect 112628 99356 112680 99408
rect 114698 99900 114750 99952
rect 114882 99900 114934 99952
rect 115158 99900 115210 99952
rect 114974 99832 115026 99884
rect 114468 99424 114520 99476
rect 115112 99628 115164 99680
rect 115020 99560 115072 99612
rect 115342 99900 115394 99952
rect 115434 99900 115486 99952
rect 115710 99764 115762 99816
rect 115480 99628 115532 99680
rect 114928 99492 114980 99544
rect 115204 99492 115256 99544
rect 115388 99492 115440 99544
rect 115664 99492 115716 99544
rect 115894 99900 115946 99952
rect 115986 99900 116038 99952
rect 116078 99900 116130 99952
rect 116262 99832 116314 99884
rect 116124 99696 116176 99748
rect 116446 99900 116498 99952
rect 116630 99900 116682 99952
rect 116722 99900 116774 99952
rect 116814 99900 116866 99952
rect 116998 99900 117050 99952
rect 116492 99764 116544 99816
rect 116584 99696 116636 99748
rect 116032 99560 116084 99612
rect 115848 99492 115900 99544
rect 115940 99492 115992 99544
rect 116308 99628 116360 99680
rect 116860 99628 116912 99680
rect 116768 99560 116820 99612
rect 117366 99900 117418 99952
rect 117458 99900 117510 99952
rect 117550 99900 117602 99952
rect 117274 99832 117326 99884
rect 117136 99628 117188 99680
rect 117826 99900 117878 99952
rect 117918 99900 117970 99952
rect 118378 99900 118430 99952
rect 118654 99900 118706 99952
rect 117504 99696 117556 99748
rect 117412 99560 117464 99612
rect 117504 99492 117556 99544
rect 117228 99424 117280 99476
rect 117320 99424 117372 99476
rect 117688 99696 117740 99748
rect 118010 99832 118062 99884
rect 118194 99832 118246 99884
rect 117872 99628 117924 99680
rect 118240 99696 118292 99748
rect 117964 99560 118016 99612
rect 118746 99832 118798 99884
rect 118424 99560 118476 99612
rect 119206 99900 119258 99952
rect 119482 99900 119534 99952
rect 119574 99900 119626 99952
rect 119666 99900 119718 99952
rect 120034 99900 120086 99952
rect 120126 99900 120178 99952
rect 120494 99900 120546 99952
rect 120586 99900 120638 99952
rect 120678 99900 120730 99952
rect 120954 99900 121006 99952
rect 118976 99560 119028 99612
rect 119850 99832 119902 99884
rect 119942 99832 119994 99884
rect 119298 99764 119350 99816
rect 119528 99764 119580 99816
rect 119620 99764 119672 99816
rect 119712 99764 119764 99816
rect 119804 99696 119856 99748
rect 119620 99628 119672 99680
rect 119896 99628 119948 99680
rect 120724 99764 120776 99816
rect 120540 99696 120592 99748
rect 120632 99696 120684 99748
rect 120816 99628 120868 99680
rect 117780 99492 117832 99544
rect 118792 99492 118844 99544
rect 120172 99560 120224 99612
rect 121598 100104 121650 100156
rect 127992 100104 128044 100156
rect 121322 100036 121374 100088
rect 125738 100036 125790 100088
rect 127118 100036 127170 100088
rect 127808 100036 127860 100088
rect 121230 99764 121282 99816
rect 121184 99628 121236 99680
rect 122794 99968 122846 100020
rect 124726 99968 124778 100020
rect 121414 99900 121466 99952
rect 121552 99628 121604 99680
rect 121460 99560 121512 99612
rect 121874 99832 121926 99884
rect 121736 99492 121788 99544
rect 122242 99900 122294 99952
rect 122334 99900 122386 99952
rect 122380 99628 122432 99680
rect 122288 99560 122340 99612
rect 122702 99900 122754 99952
rect 118332 99424 118384 99476
rect 119436 99424 119488 99476
rect 121000 99424 121052 99476
rect 122656 99492 122708 99544
rect 123254 99900 123306 99952
rect 123438 99900 123490 99952
rect 123530 99900 123582 99952
rect 123070 99832 123122 99884
rect 122932 99628 122984 99680
rect 123300 99628 123352 99680
rect 123116 99560 123168 99612
rect 123714 99832 123766 99884
rect 123576 99492 123628 99544
rect 122748 99424 122800 99476
rect 123392 99424 123444 99476
rect 123990 99900 124042 99952
rect 124082 99900 124134 99952
rect 124174 99832 124226 99884
rect 124358 99832 124410 99884
rect 124036 99696 124088 99748
rect 123852 99628 123904 99680
rect 123944 99628 123996 99680
rect 124680 99764 124732 99816
rect 124312 99696 124364 99748
rect 124404 99696 124456 99748
rect 124496 99628 124548 99680
rect 124220 99492 124272 99544
rect 125554 99900 125606 99952
rect 114744 99288 114796 99340
rect 116492 99288 116544 99340
rect 125830 99764 125882 99816
rect 126014 99900 126066 99952
rect 126290 99900 126342 99952
rect 126382 99900 126434 99952
rect 126934 99900 126986 99952
rect 127026 99900 127078 99952
rect 127210 99900 127262 99952
rect 126842 99832 126894 99884
rect 126244 99696 126296 99748
rect 125968 99560 126020 99612
rect 126244 99492 126296 99544
rect 126428 99560 126480 99612
rect 127072 99696 127124 99748
rect 127624 99832 127676 99884
rect 126888 99560 126940 99612
rect 127256 99560 127308 99612
rect 126520 99492 126572 99544
rect 125692 99356 125744 99408
rect 126152 99356 126204 99408
rect 126428 99356 126480 99408
rect 128084 99288 128136 99340
rect 116676 99084 116728 99136
rect 120080 98540 120132 98592
rect 121368 98540 121420 98592
rect 88616 98472 88668 98524
rect 88892 98472 88944 98524
rect 95240 98472 95292 98524
rect 95424 98472 95476 98524
rect 89260 98336 89312 98388
rect 90916 98336 90968 98388
rect 102048 98336 102100 98388
rect 103244 98336 103296 98388
rect 82728 98268 82780 98320
rect 86592 98268 86644 98320
rect 89720 98268 89772 98320
rect 89904 98268 89956 98320
rect 117136 98268 117188 98320
rect 117596 98268 117648 98320
rect 127348 98268 127400 98320
rect 127716 98268 127768 98320
rect 83372 98132 83424 98184
rect 83924 98132 83976 98184
rect 89444 98132 89496 98184
rect 89720 98132 89772 98184
rect 91468 98132 91520 98184
rect 90088 98064 90140 98116
rect 91744 98064 91796 98116
rect 103612 98132 103664 98184
rect 103796 98132 103848 98184
rect 110972 98064 111024 98116
rect 114284 98064 114336 98116
rect 91100 97860 91152 97912
rect 92112 97860 92164 97912
rect 92388 97860 92440 97912
rect 110972 97928 111024 97980
rect 111156 97928 111208 97980
rect 113088 97928 113140 97980
rect 113824 97928 113876 97980
rect 117964 97928 118016 97980
rect 129188 97928 129240 97980
rect 82084 97792 82136 97844
rect 98460 97792 98512 97844
rect 98828 97792 98880 97844
rect 129740 97860 129792 97912
rect 131120 97792 131172 97844
rect 81992 97724 82044 97776
rect 64880 97656 64932 97708
rect 81808 97656 81860 97708
rect 62764 97588 62816 97640
rect 84292 97588 84344 97640
rect 58624 97520 58676 97572
rect 84384 97520 84436 97572
rect 92020 97724 92072 97776
rect 92388 97724 92440 97776
rect 89996 97656 90048 97708
rect 91100 97656 91152 97708
rect 91652 97656 91704 97708
rect 131764 97724 131816 97776
rect 93584 97656 93636 97708
rect 133880 97656 133932 97708
rect 88432 97588 88484 97640
rect 89076 97588 89128 97640
rect 92204 97588 92256 97640
rect 135904 97588 135956 97640
rect 92480 97520 92532 97572
rect 92848 97520 92900 97572
rect 93492 97520 93544 97572
rect 98552 97520 98604 97572
rect 99196 97520 99248 97572
rect 104900 97520 104952 97572
rect 113824 97520 113876 97572
rect 53104 97452 53156 97504
rect 79784 97452 79836 97504
rect 85764 97452 85816 97504
rect 86132 97452 86184 97504
rect 106188 97452 106240 97504
rect 113916 97452 113968 97504
rect 54484 97384 54536 97436
rect 77852 97384 77904 97436
rect 84384 97384 84436 97436
rect 86408 97384 86460 97436
rect 90824 97384 90876 97436
rect 92020 97384 92072 97436
rect 101956 97384 102008 97436
rect 118148 97520 118200 97572
rect 121368 97520 121420 97572
rect 200764 97520 200816 97572
rect 127072 97452 127124 97504
rect 209044 97452 209096 97504
rect 118976 97384 119028 97436
rect 119344 97384 119396 97436
rect 122748 97384 122800 97436
rect 278044 97384 278096 97436
rect 43444 97316 43496 97368
rect 80428 97316 80480 97368
rect 31024 97248 31076 97300
rect 82820 97248 82872 97300
rect 93400 97248 93452 97300
rect 95056 97248 95108 97300
rect 116400 97316 116452 97368
rect 120080 97316 120132 97368
rect 120724 97316 120776 97368
rect 104900 97248 104952 97300
rect 105544 97248 105596 97300
rect 110420 97248 110472 97300
rect 81532 97180 81584 97232
rect 91008 97180 91060 97232
rect 93676 97180 93728 97232
rect 94964 97180 95016 97232
rect 89536 97112 89588 97164
rect 90456 97112 90508 97164
rect 97264 97112 97316 97164
rect 97540 97112 97592 97164
rect 81808 97044 81860 97096
rect 87788 97044 87840 97096
rect 91560 97044 91612 97096
rect 94780 97044 94832 97096
rect 71044 96976 71096 97028
rect 85488 96976 85540 97028
rect 82176 96908 82228 96960
rect 93400 96772 93452 96824
rect 82636 96636 82688 96688
rect 83096 96636 83148 96688
rect 85672 96568 85724 96620
rect 87420 96704 87472 96756
rect 86408 96636 86460 96688
rect 87512 96636 87564 96688
rect 92480 96636 92532 96688
rect 93400 96636 93452 96688
rect 110604 97112 110656 97164
rect 111156 97112 111208 97164
rect 105176 96976 105228 97028
rect 105452 96976 105504 97028
rect 118976 97248 119028 97300
rect 119620 97248 119672 97300
rect 119712 97248 119764 97300
rect 295984 97316 296036 97368
rect 124496 97248 124548 97300
rect 446404 97248 446456 97300
rect 118608 97180 118660 97232
rect 129096 97180 129148 97232
rect 119160 97112 119212 97164
rect 129280 97112 129332 97164
rect 118148 97044 118200 97096
rect 119804 97044 119856 97096
rect 121092 96976 121144 97028
rect 114928 96908 114980 96960
rect 105176 96840 105228 96892
rect 105636 96840 105688 96892
rect 118792 96908 118844 96960
rect 119160 96908 119212 96960
rect 120816 96908 120868 96960
rect 121000 96908 121052 96960
rect 118884 96840 118936 96892
rect 119528 96840 119580 96892
rect 111616 96772 111668 96824
rect 112812 96772 112864 96824
rect 113088 96772 113140 96824
rect 114928 96772 114980 96824
rect 115756 96772 115808 96824
rect 117044 96772 117096 96824
rect 118516 96772 118568 96824
rect 118792 96772 118844 96824
rect 119436 96772 119488 96824
rect 106464 96704 106516 96756
rect 107108 96704 107160 96756
rect 113824 96704 113876 96756
rect 119712 96704 119764 96756
rect 120356 96704 120408 96756
rect 127992 96704 128044 96756
rect 121368 96636 121420 96688
rect 123576 96636 123628 96688
rect 125140 96636 125192 96688
rect 82268 96500 82320 96552
rect 95332 96568 95384 96620
rect 106280 96568 106332 96620
rect 106740 96568 106792 96620
rect 109132 96568 109184 96620
rect 110236 96568 110288 96620
rect 118884 96568 118936 96620
rect 119620 96568 119672 96620
rect 103520 96500 103572 96552
rect 103888 96500 103940 96552
rect 116400 96500 116452 96552
rect 116860 96500 116912 96552
rect 117688 96500 117740 96552
rect 127900 96500 127952 96552
rect 94872 96432 94924 96484
rect 129004 96568 129056 96620
rect 81348 96364 81400 96416
rect 94228 96364 94280 96416
rect 94688 96364 94740 96416
rect 101036 96364 101088 96416
rect 135996 96364 136048 96416
rect 80980 96296 81032 96348
rect 93768 96296 93820 96348
rect 94596 96296 94648 96348
rect 95240 96296 95292 96348
rect 176660 96296 176712 96348
rect 81440 96228 81492 96280
rect 96436 96228 96488 96280
rect 96620 96228 96672 96280
rect 193220 96228 193272 96280
rect 82360 96160 82412 96212
rect 95976 96160 96028 96212
rect 97448 96160 97500 96212
rect 200120 96160 200172 96212
rect 106832 96092 106884 96144
rect 81256 96024 81308 96076
rect 93216 96024 93268 96076
rect 103520 96024 103572 96076
rect 103704 96024 103756 96076
rect 106372 96024 106424 96076
rect 107016 96024 107068 96076
rect 105084 95956 105136 96008
rect 105728 95956 105780 96008
rect 106280 95956 106332 96008
rect 106832 95956 106884 96008
rect 107016 95888 107068 95940
rect 107384 96092 107436 96144
rect 107936 96092 107988 96144
rect 109040 96092 109092 96144
rect 109500 96092 109552 96144
rect 114928 96092 114980 96144
rect 115756 96092 115808 96144
rect 117504 96092 117556 96144
rect 117688 96092 117740 96144
rect 122012 96092 122064 96144
rect 498200 96092 498252 96144
rect 109224 96024 109276 96076
rect 109868 96024 109920 96076
rect 123852 96024 123904 96076
rect 514760 96024 514812 96076
rect 114928 95956 114980 96008
rect 115112 95956 115164 96008
rect 125508 95956 125560 96008
rect 528560 95956 528612 96008
rect 126520 95888 126572 95940
rect 545120 95888 545172 95940
rect 81164 95820 81216 95872
rect 93308 95820 93360 95872
rect 96712 95820 96764 95872
rect 97172 95820 97224 95872
rect 105084 95820 105136 95872
rect 105360 95820 105412 95872
rect 106280 95820 106332 95872
rect 107200 95820 107252 95872
rect 81072 95752 81124 95804
rect 93584 95752 93636 95804
rect 94504 95752 94556 95804
rect 103612 95752 103664 95804
rect 104348 95752 104400 95804
rect 116952 95752 117004 95804
rect 122472 95752 122524 95804
rect 104992 95684 105044 95736
rect 105360 95684 105412 95736
rect 109408 95616 109460 95668
rect 109960 95616 110012 95668
rect 102140 95548 102192 95600
rect 102600 95548 102652 95600
rect 104992 95548 105044 95600
rect 105176 95548 105228 95600
rect 107752 95548 107804 95600
rect 108764 95548 108816 95600
rect 110512 95548 110564 95600
rect 111524 95548 111576 95600
rect 102232 95412 102284 95464
rect 102600 95412 102652 95464
rect 115848 95344 115900 95396
rect 118148 95344 118200 95396
rect 121552 95344 121604 95396
rect 121920 95344 121972 95396
rect 95332 95208 95384 95260
rect 96160 95208 96212 95260
rect 114836 95140 114888 95192
rect 115480 95140 115532 95192
rect 121460 95140 121512 95192
rect 121828 95140 121880 95192
rect 110236 95072 110288 95124
rect 115848 95072 115900 95124
rect 113456 95004 113508 95056
rect 113824 95004 113876 95056
rect 116032 95004 116084 95056
rect 116400 95004 116452 95056
rect 91284 94936 91336 94988
rect 126980 95004 127032 95056
rect 121644 94936 121696 94988
rect 122564 94936 122616 94988
rect 123300 94936 123352 94988
rect 123484 94936 123536 94988
rect 107476 94868 107528 94920
rect 162124 94868 162176 94920
rect 96620 94800 96672 94852
rect 97908 94800 97960 94852
rect 101220 94800 101272 94852
rect 247040 94800 247092 94852
rect 84752 94732 84804 94784
rect 85120 94732 85172 94784
rect 88708 94732 88760 94784
rect 89076 94732 89128 94784
rect 101864 94732 101916 94784
rect 252560 94732 252612 94784
rect 81532 94664 81584 94716
rect 82452 94664 82504 94716
rect 83372 94664 83424 94716
rect 83648 94664 83700 94716
rect 85028 94664 85080 94716
rect 85396 94664 85448 94716
rect 87144 94664 87196 94716
rect 87236 94664 87288 94716
rect 87512 94664 87564 94716
rect 88800 94664 88852 94716
rect 95884 94664 95936 94716
rect 96344 94664 96396 94716
rect 96804 94664 96856 94716
rect 98092 94664 98144 94716
rect 99288 94664 99340 94716
rect 103336 94664 103388 94716
rect 266360 94664 266412 94716
rect 83096 94528 83148 94580
rect 83464 94528 83516 94580
rect 85856 94528 85908 94580
rect 86316 94528 86368 94580
rect 86960 94528 87012 94580
rect 87604 94528 87656 94580
rect 87420 94460 87472 94512
rect 88064 94460 88116 94512
rect 82912 94392 82964 94444
rect 83464 94392 83516 94444
rect 83556 94392 83608 94444
rect 83740 94392 83792 94444
rect 84844 94392 84896 94444
rect 85304 94392 85356 94444
rect 85856 94392 85908 94444
rect 86868 94392 86920 94444
rect 87144 94392 87196 94444
rect 87880 94392 87932 94444
rect 84384 94324 84436 94376
rect 84936 94324 84988 94376
rect 85948 94324 86000 94376
rect 86776 94324 86828 94376
rect 88064 94324 88116 94376
rect 88340 94528 88392 94580
rect 88340 94392 88392 94444
rect 91376 94596 91428 94648
rect 91836 94596 91888 94648
rect 90088 94528 90140 94580
rect 90272 94528 90324 94580
rect 91284 94528 91336 94580
rect 91928 94528 91980 94580
rect 93860 94528 93912 94580
rect 94044 94528 94096 94580
rect 94228 94528 94280 94580
rect 94412 94528 94464 94580
rect 95516 94528 95568 94580
rect 95792 94528 95844 94580
rect 95884 94528 95936 94580
rect 96068 94528 96120 94580
rect 98000 94596 98052 94648
rect 98368 94596 98420 94648
rect 106004 94596 106056 94648
rect 296720 94596 296772 94648
rect 98092 94528 98144 94580
rect 98276 94528 98328 94580
rect 100024 94528 100076 94580
rect 100668 94528 100720 94580
rect 100944 94528 100996 94580
rect 101588 94528 101640 94580
rect 109592 94528 109644 94580
rect 111800 94528 111852 94580
rect 111984 94528 112036 94580
rect 112076 94528 112128 94580
rect 89904 94460 89956 94512
rect 90640 94460 90692 94512
rect 91836 94460 91888 94512
rect 92388 94460 92440 94512
rect 96804 94460 96856 94512
rect 96896 94460 96948 94512
rect 97356 94460 97408 94512
rect 108948 94460 109000 94512
rect 89812 94392 89864 94444
rect 90272 94392 90324 94444
rect 91100 94392 91152 94444
rect 91928 94392 91980 94444
rect 93768 94392 93820 94444
rect 94044 94392 94096 94444
rect 101036 94392 101088 94444
rect 101220 94392 101272 94444
rect 108856 94392 108908 94444
rect 109592 94392 109644 94444
rect 88524 94324 88576 94376
rect 88616 94324 88668 94376
rect 89628 94324 89680 94376
rect 92572 94324 92624 94376
rect 93032 94324 93084 94376
rect 95976 94324 96028 94376
rect 96528 94324 96580 94376
rect 98368 94324 98420 94376
rect 98736 94324 98788 94376
rect 112168 94324 112220 94376
rect 112536 94324 112588 94376
rect 89812 94256 89864 94308
rect 90548 94256 90600 94308
rect 97908 94256 97960 94308
rect 98460 94256 98512 94308
rect 112076 94256 112128 94308
rect 112444 94256 112496 94308
rect 92572 94188 92624 94240
rect 93676 94188 93728 94240
rect 112536 94188 112588 94240
rect 116032 94528 116084 94580
rect 116308 94528 116360 94580
rect 113548 94460 113600 94512
rect 113732 94460 113784 94512
rect 115204 94460 115256 94512
rect 115388 94460 115440 94512
rect 115848 94460 115900 94512
rect 342260 94528 342312 94580
rect 113272 94392 113324 94444
rect 114100 94392 114152 94444
rect 114560 94392 114612 94444
rect 115112 94392 115164 94444
rect 116308 94392 116360 94444
rect 116768 94392 116820 94444
rect 118332 94392 118384 94444
rect 118516 94392 118568 94444
rect 113088 94324 113140 94376
rect 113732 94324 113784 94376
rect 114744 94324 114796 94376
rect 115572 94324 115624 94376
rect 117320 94324 117372 94376
rect 117872 94324 117924 94376
rect 114468 94256 114520 94308
rect 398840 94460 398892 94512
rect 121920 94392 121972 94444
rect 122288 94392 122340 94444
rect 122932 94392 122984 94444
rect 123300 94392 123352 94444
rect 124496 94392 124548 94444
rect 124772 94392 124824 94444
rect 123024 94324 123076 94376
rect 123392 94324 123444 94376
rect 121644 94256 121696 94308
rect 122380 94256 122432 94308
rect 122748 94256 122800 94308
rect 123300 94256 123352 94308
rect 124404 94256 124456 94308
rect 124772 94256 124824 94308
rect 123024 94188 123076 94240
rect 123760 94188 123812 94240
rect 107844 94120 107896 94172
rect 108488 94120 108540 94172
rect 111708 94120 111760 94172
rect 112444 94120 112496 94172
rect 120172 94120 120224 94172
rect 121276 94120 121328 94172
rect 124404 94120 124456 94172
rect 125048 94120 125100 94172
rect 107844 93984 107896 94036
rect 108212 93984 108264 94036
rect 105176 93916 105228 93968
rect 105912 93916 105964 93968
rect 119528 93780 119580 93832
rect 128084 93780 128136 93832
rect 110328 93712 110380 93764
rect 111524 93712 111576 93764
rect 108028 93440 108080 93492
rect 329840 93440 329892 93492
rect 111340 93372 111392 93424
rect 346400 93372 346452 93424
rect 109776 93304 109828 93356
rect 349160 93304 349212 93356
rect 112812 93236 112864 93288
rect 374000 93236 374052 93288
rect 114376 93168 114428 93220
rect 391940 93168 391992 93220
rect 115756 93100 115808 93152
rect 401600 93100 401652 93152
rect 103428 92760 103480 92812
rect 104256 92760 104308 92812
rect 101036 92488 101088 92540
rect 101680 92488 101732 92540
rect 97264 92420 97316 92472
rect 128820 92420 128872 92472
rect 93400 92352 93452 92404
rect 142160 92352 142212 92404
rect 121368 92284 121420 92336
rect 171140 92284 171192 92336
rect 116860 92216 116912 92268
rect 175280 92216 175332 92268
rect 97172 92148 97224 92200
rect 125048 92148 125100 92200
rect 128820 92148 128872 92200
rect 194600 92148 194652 92200
rect 99472 92080 99524 92132
rect 128912 92080 128964 92132
rect 224960 92080 225012 92132
rect 121092 92012 121144 92064
rect 357440 92012 357492 92064
rect 114284 91944 114336 91996
rect 362960 91944 363012 91996
rect 118608 91876 118660 91928
rect 445760 91876 445812 91928
rect 119344 91808 119396 91860
rect 456800 91808 456852 91860
rect 90364 91740 90416 91792
rect 120264 91740 120316 91792
rect 125140 91740 125192 91792
rect 506480 91740 506532 91792
rect 125048 91060 125100 91112
rect 191840 91060 191892 91112
rect 98828 90992 98880 91044
rect 128728 90992 128780 91044
rect 94596 90652 94648 90704
rect 158720 90652 158772 90704
rect 128728 90584 128780 90636
rect 211160 90584 211212 90636
rect 119712 90516 119764 90568
rect 291200 90516 291252 90568
rect 113916 90448 113968 90500
rect 307760 90448 307812 90500
rect 107108 90380 107160 90432
rect 310520 90380 310572 90432
rect 91468 90312 91520 90364
rect 119344 90312 119396 90364
rect 120908 90312 120960 90364
rect 473452 90312 473504 90364
rect 107936 90244 107988 90296
rect 108304 90244 108356 90296
rect 108028 90176 108080 90228
rect 108580 90176 108632 90228
rect 102416 90108 102468 90160
rect 102968 90108 103020 90160
rect 108304 90108 108356 90160
rect 108488 90108 108540 90160
rect 114560 89972 114612 90024
rect 115664 89972 115716 90024
rect 98552 89632 98604 89684
rect 128360 89632 128412 89684
rect 92572 89564 92624 89616
rect 144920 89564 144972 89616
rect 96160 89496 96212 89548
rect 178040 89496 178092 89548
rect 95884 89428 95936 89480
rect 180800 89428 180852 89480
rect 128360 89360 128412 89412
rect 128636 89360 128688 89412
rect 218060 89360 218112 89412
rect 119804 89292 119856 89344
rect 129832 89292 129884 89344
rect 241520 89292 241572 89344
rect 103244 89224 103296 89276
rect 258080 89224 258132 89276
rect 104532 89156 104584 89208
rect 287060 89156 287112 89208
rect 105728 89088 105780 89140
rect 293960 89088 294012 89140
rect 115388 89020 115440 89072
rect 409880 89020 409932 89072
rect 116676 88952 116728 89004
rect 429200 88952 429252 89004
rect 127256 88884 127308 88936
rect 127532 88884 127584 88936
rect 98460 88272 98512 88324
rect 128452 88272 128504 88324
rect 208400 88272 208452 88324
rect 99932 88204 99984 88256
rect 128544 88204 128596 88256
rect 227720 88204 227772 88256
rect 101496 88136 101548 88188
rect 251180 88136 251232 88188
rect 111156 88068 111208 88120
rect 360200 88068 360252 88120
rect 200764 88000 200816 88052
rect 469220 88000 469272 88052
rect 115296 87932 115348 87984
rect 407120 87932 407172 87984
rect 118424 87864 118476 87916
rect 429292 87864 429344 87916
rect 123576 87796 123628 87848
rect 512000 87796 512052 87848
rect 77300 87728 77352 87780
rect 88064 87728 88116 87780
rect 123668 87728 123720 87780
rect 516140 87728 516192 87780
rect 56600 87660 56652 87712
rect 85488 87660 85540 87712
rect 126428 87660 126480 87712
rect 545212 87660 545264 87712
rect 40040 87592 40092 87644
rect 84016 87592 84068 87644
rect 91376 87592 91428 87644
rect 115388 87592 115440 87644
rect 126336 87592 126388 87644
rect 549260 87592 549312 87644
rect 101404 86572 101456 86624
rect 244280 86572 244332 86624
rect 101312 86504 101364 86556
rect 247132 86504 247184 86556
rect 104256 86436 104308 86488
rect 274640 86436 274692 86488
rect 104348 86368 104400 86420
rect 282920 86368 282972 86420
rect 116584 86300 116636 86352
rect 433340 86300 433392 86352
rect 53840 86232 53892 86284
rect 85212 86232 85264 86284
rect 117780 86232 117832 86284
rect 445852 86232 445904 86284
rect 97080 85484 97132 85536
rect 128360 85484 128412 85536
rect 197360 85212 197412 85264
rect 94320 85144 94372 85196
rect 164240 85144 164292 85196
rect 108764 85076 108816 85128
rect 324320 85076 324372 85128
rect 112536 85008 112588 85060
rect 376760 85008 376812 85060
rect 112628 84940 112680 84992
rect 379520 84940 379572 84992
rect 31760 84872 31812 84924
rect 83924 84872 83976 84924
rect 116492 84872 116544 84924
rect 426440 84872 426492 84924
rect 117688 84804 117740 84856
rect 440240 84804 440292 84856
rect 83556 84192 83608 84244
rect 86408 84192 86460 84244
rect 75920 83444 75972 83496
rect 85580 83444 85632 83496
rect 109684 83444 109736 83496
rect 345020 83444 345072 83496
rect 100300 82288 100352 82340
rect 100576 82288 100628 82340
rect 107016 82220 107068 82272
rect 313280 82220 313332 82272
rect 113824 82152 113876 82204
rect 390560 82152 390612 82204
rect 123484 82084 123536 82136
rect 512092 82084 512144 82136
rect 122472 80724 122524 80776
rect 434720 80724 434772 80776
rect 123392 80656 123444 80708
rect 507860 80656 507912 80708
rect 136088 71680 136140 71732
rect 579620 71680 579672 71732
rect 129280 54476 129332 54528
rect 462320 54476 462372 54528
rect 129188 53116 129240 53168
rect 448520 53116 448572 53168
rect 129096 53048 129148 53100
rect 455420 53048 455472 53100
rect 89168 46248 89220 46300
rect 100024 46248 100076 46300
rect 99840 46180 99892 46232
rect 225052 46180 225104 46232
rect 70400 44956 70452 45008
rect 82636 44956 82688 45008
rect 46940 44888 46992 44940
rect 84752 44888 84804 44940
rect 30380 44820 30432 44872
rect 82544 44820 82596 44872
rect 94780 42100 94832 42152
rect 131212 42100 131264 42152
rect 91284 42032 91336 42084
rect 136732 42032 136784 42084
rect 94228 41148 94280 41200
rect 165620 41148 165672 41200
rect 101220 41080 101272 41132
rect 242900 41080 242952 41132
rect 105636 41012 105688 41064
rect 302240 41012 302292 41064
rect 105544 40944 105596 40996
rect 302332 40944 302384 40996
rect 116400 40876 116452 40928
rect 423680 40876 423732 40928
rect 119160 40808 119212 40860
rect 456892 40808 456944 40860
rect 119068 40740 119120 40792
rect 460940 40740 460992 40792
rect 119252 40672 119304 40724
rect 465080 40672 465132 40724
rect 100484 39720 100536 39772
rect 237380 39720 237432 39772
rect 109592 39652 109644 39704
rect 340880 39652 340932 39704
rect 112444 39584 112496 39636
rect 374092 39584 374144 39636
rect 117596 39516 117648 39568
rect 443000 39516 443052 39568
rect 120816 39448 120868 39500
rect 483020 39448 483072 39500
rect 124956 39380 125008 39432
rect 532700 39380 532752 39432
rect 126244 39312 126296 39364
rect 542360 39312 542412 39364
rect 99656 38224 99708 38276
rect 230480 38224 230532 38276
rect 99748 38156 99800 38208
rect 233240 38156 233292 38208
rect 118332 38088 118384 38140
rect 415400 38088 415452 38140
rect 116952 38020 117004 38072
rect 422300 38020 422352 38072
rect 116216 37952 116268 38004
rect 425060 37952 425112 38004
rect 116308 37884 116360 37936
rect 431960 37884 432012 37936
rect 95700 36660 95752 36712
rect 180892 36660 180944 36712
rect 96988 36592 97040 36644
rect 197452 36592 197504 36644
rect 118240 36524 118292 36576
rect 408500 36524 408552 36576
rect 115204 35436 115256 35488
rect 418160 35436 418212 35488
rect 117504 35368 117556 35420
rect 440332 35368 440384 35420
rect 117412 35300 117464 35352
rect 444380 35300 444432 35352
rect 120724 35232 120776 35284
rect 478880 35232 478932 35284
rect 124864 35164 124916 35216
rect 531320 35164 531372 35216
rect 111064 34280 111116 34332
rect 363052 34280 363104 34332
rect 110972 34212 111024 34264
rect 365720 34212 365772 34264
rect 115112 34144 115164 34196
rect 407212 34144 407264 34196
rect 115020 34076 115072 34128
rect 411260 34076 411312 34128
rect 114928 34008 114980 34060
rect 414020 34008 414072 34060
rect 116032 33940 116084 33992
rect 427820 33940 427872 33992
rect 116124 33872 116176 33924
rect 430580 33872 430632 33924
rect 117320 33804 117372 33856
rect 447140 33804 447192 33856
rect 120632 33736 120684 33788
rect 481640 33736 481692 33788
rect 98368 32852 98420 32904
rect 216680 32852 216732 32904
rect 108396 32784 108448 32836
rect 332600 32784 332652 32836
rect 112260 32716 112312 32768
rect 378140 32716 378192 32768
rect 112352 32648 112404 32700
rect 380900 32648 380952 32700
rect 112168 32580 112220 32632
rect 385132 32580 385184 32632
rect 113732 32512 113784 32564
rect 390652 32512 390704 32564
rect 113640 32444 113692 32496
rect 394700 32444 394752 32496
rect 113548 32376 113600 32428
rect 397460 32376 397512 32428
rect 94044 31492 94096 31544
rect 158812 31492 158864 31544
rect 94136 31424 94188 31476
rect 162860 31424 162912 31476
rect 106924 31356 106976 31408
rect 316040 31356 316092 31408
rect 108304 31288 108356 31340
rect 325700 31288 325752 31340
rect 109500 31220 109552 31272
rect 340972 31220 341024 31272
rect 111432 31152 111484 31204
rect 354680 31152 354732 31204
rect 110788 31084 110840 31136
rect 361580 31084 361632 31136
rect 110880 31016 110932 31068
rect 364340 31016 364392 31068
rect 93952 30132 94004 30184
rect 160100 30132 160152 30184
rect 106740 30064 106792 30116
rect 307852 30064 307904 30116
rect 106832 29996 106884 30048
rect 309140 29996 309192 30048
rect 106556 29928 106608 29980
rect 311900 29928 311952 29980
rect 106648 29860 106700 29912
rect 313372 29860 313424 29912
rect 106464 29792 106516 29844
rect 314660 29792 314712 29844
rect 108120 29724 108172 29776
rect 324412 29724 324464 29776
rect 108212 29656 108264 29708
rect 328460 29656 328512 29708
rect 120540 29588 120592 29640
rect 478972 29588 479024 29640
rect 104072 28636 104124 28688
rect 276020 28636 276072 28688
rect 103980 28568 104032 28620
rect 280160 28568 280212 28620
rect 104164 28500 104216 28552
rect 281540 28500 281592 28552
rect 105360 28432 105412 28484
rect 291292 28432 291344 28484
rect 105452 28364 105504 28416
rect 295340 28364 295392 28416
rect 105268 28296 105320 28348
rect 299480 28296 299532 28348
rect 110696 28228 110748 28280
rect 357532 28228 357584 28280
rect 92848 27276 92900 27328
rect 149060 27276 149112 27328
rect 92940 27208 92992 27260
rect 150440 27208 150492 27260
rect 102876 27140 102928 27192
rect 258172 27140 258224 27192
rect 102692 27072 102744 27124
rect 262220 27072 262272 27124
rect 102784 27004 102836 27056
rect 264980 27004 265032 27056
rect 103888 26936 103940 26988
rect 274732 26936 274784 26988
rect 103796 26868 103848 26920
rect 278780 26868 278832 26920
rect 92756 26052 92808 26104
rect 146300 26052 146352 26104
rect 100852 25984 100904 26036
rect 241612 25984 241664 26036
rect 101128 25916 101180 25968
rect 245660 25916 245712 25968
rect 100944 25848 100996 25900
rect 248420 25848 248472 25900
rect 101036 25780 101088 25832
rect 252652 25780 252704 25832
rect 111892 25712 111944 25764
rect 375380 25712 375432 25764
rect 111984 25644 112036 25696
rect 379612 25644 379664 25696
rect 112076 25576 112128 25628
rect 382280 25576 382332 25628
rect 113456 25508 113508 25560
rect 396080 25508 396132 25560
rect 92664 24488 92716 24540
rect 142252 24488 142304 24540
rect 96896 24420 96948 24472
rect 198740 24420 198792 24472
rect 98184 24352 98236 24404
rect 208492 24352 208544 24404
rect 98092 24284 98144 24336
rect 212540 24284 212592 24336
rect 98276 24216 98328 24268
rect 215300 24216 215352 24268
rect 110604 24148 110656 24200
rect 358820 24148 358872 24200
rect 118976 24080 119028 24132
rect 463700 24080 463752 24132
rect 95608 23128 95660 23180
rect 179420 23128 179472 23180
rect 95516 23060 95568 23112
rect 182180 23060 182232 23112
rect 96804 22992 96856 23044
rect 191932 22992 191984 23044
rect 96712 22924 96764 22976
rect 195980 22924 196032 22976
rect 100760 22856 100812 22908
rect 249800 22856 249852 22908
rect 102600 22788 102652 22840
rect 259460 22788 259512 22840
rect 102508 22720 102560 22772
rect 263600 22720 263652 22772
rect 93584 21836 93636 21888
rect 147680 21836 147732 21888
rect 95424 21768 95476 21820
rect 175372 21768 175424 21820
rect 99564 21700 99616 21752
rect 226340 21700 226392 21752
rect 123300 21632 123352 21684
rect 506572 21632 506624 21684
rect 123208 21564 123260 21616
rect 510620 21564 510672 21616
rect 123116 21496 123168 21548
rect 513380 21496 513432 21548
rect 124772 21428 124824 21480
rect 523132 21428 523184 21480
rect 38660 21360 38712 21412
rect 83648 21360 83700 21412
rect 90272 21360 90324 21412
rect 110604 21360 110656 21412
rect 126152 21360 126204 21412
rect 550640 21360 550692 21412
rect 98000 20408 98052 20460
rect 213920 20408 213972 20460
rect 122104 20340 122156 20392
rect 490012 20340 490064 20392
rect 122012 20272 122064 20324
rect 494060 20272 494112 20324
rect 122196 20204 122248 20256
rect 496820 20204 496872 20256
rect 121920 20136 121972 20188
rect 500960 20136 501012 20188
rect 126060 20068 126112 20120
rect 546500 20068 546552 20120
rect 84752 20000 84804 20052
rect 87788 20000 87840 20052
rect 127808 20000 127860 20052
rect 557540 20000 557592 20052
rect 89076 19932 89128 19984
rect 98092 19932 98144 19984
rect 127440 19932 127492 19984
rect 561680 19932 561732 19984
rect 114836 18980 114888 19032
rect 169024 18980 169076 19032
rect 93860 18912 93912 18964
rect 168380 18912 168432 18964
rect 96344 18844 96396 18896
rect 183560 18844 183612 18896
rect 118884 18776 118936 18828
rect 466460 18776 466512 18828
rect 120448 18708 120500 18760
rect 477500 18708 477552 18760
rect 123024 18640 123076 18692
rect 517520 18640 517572 18692
rect 124680 18572 124732 18624
rect 524420 18572 524472 18624
rect 93032 17620 93084 17672
rect 143540 17620 143592 17672
rect 94688 17552 94740 17604
rect 164332 17552 164384 17604
rect 118700 17484 118752 17536
rect 459560 17484 459612 17536
rect 118792 17416 118844 17468
rect 462412 17416 462464 17468
rect 120356 17348 120408 17400
rect 474740 17348 474792 17400
rect 121828 17280 121880 17332
rect 491300 17280 491352 17332
rect 121736 17212 121788 17264
rect 495532 17212 495584 17264
rect 94596 16260 94648 16312
rect 162032 16260 162084 16312
rect 114652 16192 114704 16244
rect 412732 16192 412784 16244
rect 114744 16124 114796 16176
rect 417240 16124 417292 16176
rect 114560 16056 114612 16108
rect 418344 16056 418396 16108
rect 115940 15988 115992 16040
rect 423772 15988 423824 16040
rect 125968 15920 126020 15972
rect 541992 15920 542044 15972
rect 127716 15852 127768 15904
rect 560760 15852 560812 15904
rect 109408 14764 109460 14816
rect 352104 14764 352156 14816
rect 110512 14696 110564 14748
rect 368664 14696 368716 14748
rect 111800 14628 111852 14680
rect 384120 14628 384172 14680
rect 113364 14560 113416 14612
rect 394056 14560 394108 14612
rect 113180 14492 113232 14544
rect 396172 14492 396224 14544
rect 113272 14424 113324 14476
rect 400680 14424 400732 14476
rect 93308 13472 93360 13524
rect 155592 13472 155644 13524
rect 107936 13404 107988 13456
rect 332232 13404 332284 13456
rect 108028 13336 108080 13388
rect 335544 13336 335596 13388
rect 109132 13268 109184 13320
rect 344376 13268 344428 13320
rect 109316 13200 109368 13252
rect 346492 13200 346544 13252
rect 109224 13132 109276 13184
rect 351000 13132 351052 13184
rect 110420 13064 110472 13116
rect 367560 13064 367612 13116
rect 93216 12180 93268 12232
rect 152280 12180 152332 12232
rect 106372 12112 106424 12164
rect 317880 12112 317932 12164
rect 106280 12044 106332 12096
rect 318984 12044 319036 12096
rect 107660 11976 107712 12028
rect 327816 11976 327868 12028
rect 107844 11908 107896 11960
rect 329932 11908 329984 11960
rect 107752 11840 107804 11892
rect 334440 11840 334492 11892
rect 109040 11772 109092 11824
rect 348792 11772 348844 11824
rect 125876 11704 125928 11756
rect 544200 11704 544252 11756
rect 93124 10752 93176 10804
rect 147772 10752 147824 10804
rect 102416 10684 102468 10736
rect 269304 10684 269356 10736
rect 103704 10616 103756 10668
rect 280252 10616 280304 10668
rect 103612 10548 103664 10600
rect 284760 10548 284812 10600
rect 105084 10480 105136 10532
rect 296812 10480 296864 10532
rect 104992 10412 105044 10464
rect 301320 10412 301372 10464
rect 105176 10344 105228 10396
rect 304632 10344 304684 10396
rect 125784 10276 125836 10328
rect 539600 10276 539652 10328
rect 100576 9256 100628 9308
rect 235080 9256 235132 9308
rect 102324 9188 102376 9240
rect 261576 9188 261628 9240
rect 102140 9120 102192 9172
rect 264888 9120 264940 9172
rect 102232 9052 102284 9104
rect 268200 9052 268252 9104
rect 103520 8984 103572 9036
rect 278136 8984 278188 9036
rect 209044 8916 209096 8968
rect 557448 8916 557500 8968
rect 97540 8100 97592 8152
rect 201960 8100 202012 8152
rect 96620 8032 96672 8084
rect 205272 8032 205324 8084
rect 98828 7964 98880 8016
rect 215208 7964 215260 8016
rect 99288 7896 99340 7948
rect 221832 7896 221884 7948
rect 99472 7828 99524 7880
rect 229560 7828 229612 7880
rect 100668 7760 100720 7812
rect 231768 7760 231820 7812
rect 124588 7692 124640 7744
rect 527640 7692 527692 7744
rect 61752 7624 61804 7676
rect 86316 7624 86368 7676
rect 124496 7624 124548 7676
rect 530952 7624 531004 7676
rect 26424 7556 26476 7608
rect 83464 7556 83516 7608
rect 124404 7556 124456 7608
rect 534264 7556 534316 7608
rect 517520 7488 517572 7540
rect 518808 7488 518860 7540
rect 523132 7488 523184 7540
rect 524328 7488 524380 7540
rect 73896 6740 73948 6792
rect 85948 6740 86000 6792
rect 70584 6672 70636 6724
rect 84936 6672 84988 6724
rect 68376 6604 68428 6656
rect 86040 6604 86092 6656
rect 67272 6536 67324 6588
rect 86224 6536 86276 6588
rect 91192 6536 91244 6588
rect 129096 6536 129148 6588
rect 63960 6468 64012 6520
rect 86132 6468 86184 6520
rect 96068 6468 96120 6520
rect 185400 6468 185452 6520
rect 62856 6400 62908 6452
rect 84844 6400 84896 6452
rect 95976 6400 96028 6452
rect 188712 6400 188764 6452
rect 55128 6332 55180 6384
rect 84660 6332 84712 6384
rect 91836 6332 91888 6384
rect 106188 6332 106240 6384
rect 122932 6332 122984 6384
rect 517704 6332 517756 6384
rect 48504 6264 48556 6316
rect 84568 6264 84620 6316
rect 91744 6264 91796 6316
rect 114744 6264 114796 6316
rect 125692 6264 125744 6316
rect 539784 6264 539836 6316
rect 38568 6196 38620 6248
rect 83372 6196 83424 6248
rect 90180 6196 90232 6248
rect 113640 6196 113692 6248
rect 127624 6196 127676 6248
rect 556344 6196 556396 6248
rect 34152 6128 34204 6180
rect 83280 6128 83332 6180
rect 90088 6128 90140 6180
rect 116952 6128 117004 6180
rect 127532 6128 127584 6180
rect 559656 6128 559708 6180
rect 88984 5448 89036 5500
rect 100392 5448 100444 5500
rect 96252 5380 96304 5432
rect 75000 5312 75052 5364
rect 85856 5312 85908 5364
rect 90824 5312 90876 5364
rect 80060 5244 80112 5296
rect 83188 5244 83240 5296
rect 88892 5244 88944 5296
rect 97080 5244 97132 5296
rect 56232 5176 56284 5228
rect 85028 5176 85080 5228
rect 89720 5176 89772 5228
rect 186504 5312 186556 5364
rect 100116 5244 100168 5296
rect 232872 5244 232924 5296
rect 52920 5108 52972 5160
rect 85396 5108 85448 5160
rect 90456 5108 90508 5160
rect 103704 5176 103756 5228
rect 104900 5176 104952 5228
rect 299112 5176 299164 5228
rect 50712 5040 50764 5092
rect 85120 5040 85172 5092
rect 89996 5040 90048 5092
rect 120172 5108 120224 5160
rect 481272 5108 481324 5160
rect 49608 4972 49660 5024
rect 84476 4972 84528 5024
rect 25320 4904 25372 4956
rect 82452 4904 82504 4956
rect 107016 5040 107068 5092
rect 121644 5040 121696 5092
rect 500040 5040 500092 5092
rect 108120 4972 108172 5024
rect 122840 4972 122892 5024
rect 509976 4972 510028 5024
rect 110328 4904 110380 4956
rect 124312 4904 124364 4956
rect 526536 4904 526588 4956
rect 24216 4836 24268 4888
rect 81624 4836 81676 4888
rect 92020 4836 92072 4888
rect 119160 4836 119212 4888
rect 124220 4836 124272 4888
rect 516784 4836 516836 4888
rect 23112 4768 23164 4820
rect 81532 4768 81584 4820
rect 82360 4768 82412 4820
rect 87696 4768 87748 4820
rect 89904 4768 89956 4820
rect 120264 4768 120316 4820
rect 125600 4768 125652 4820
rect 548616 4768 548668 4820
rect 516784 4700 516836 4752
rect 529848 4700 529900 4752
rect 88708 4292 88760 4344
rect 94872 4292 94924 4344
rect 88800 4156 88852 4208
rect 93768 4156 93820 4208
rect 75736 4088 75788 4140
rect 83740 4088 83792 4140
rect 88432 4088 88484 4140
rect 95976 4088 96028 4140
rect 131212 4088 131264 4140
rect 132408 4088 132460 4140
rect 162124 4088 162176 4140
rect 79416 4020 79468 4072
rect 87512 4020 87564 4072
rect 98644 4020 98696 4072
rect 170956 4020 171008 4072
rect 51816 3952 51868 4004
rect 62764 3952 62816 4004
rect 76104 3952 76156 4004
rect 87604 3952 87656 4004
rect 106188 3952 106240 4004
rect 139032 3952 139084 4004
rect 142252 3952 142304 4004
rect 143448 3952 143500 4004
rect 147772 3952 147824 4004
rect 148968 3952 149020 4004
rect 158812 3952 158864 4004
rect 160008 3952 160060 4004
rect 175372 4020 175424 4072
rect 176568 4020 176620 4072
rect 191932 4020 191984 4072
rect 193128 4020 193180 4072
rect 208492 4020 208544 4072
rect 209688 4020 209740 4072
rect 293592 4020 293644 4072
rect 296812 4020 296864 4072
rect 298008 4020 298060 4072
rect 307852 4020 307904 4072
rect 309048 4020 309100 4072
rect 324412 4020 324464 4072
rect 325608 4020 325660 4072
rect 329932 4020 329984 4072
rect 331128 4020 331180 4072
rect 340972 4020 341024 4072
rect 342168 4020 342220 4072
rect 346492 4020 346544 4072
rect 347688 4020 347740 4072
rect 357532 4020 357584 4072
rect 358728 4020 358780 4072
rect 390652 4020 390704 4072
rect 391848 4020 391900 4072
rect 396172 4020 396224 4072
rect 397368 4020 397420 4072
rect 407212 4020 407264 4072
rect 408408 4020 408460 4072
rect 44088 3884 44140 3936
rect 54484 3884 54536 3936
rect 58440 3884 58492 3936
rect 71044 3884 71096 3936
rect 72792 3884 72844 3936
rect 86684 3884 86736 3936
rect 94504 3884 94556 3936
rect 104808 3884 104860 3936
rect 115388 3884 115440 3936
rect 135720 3884 135772 3936
rect 135996 3884 136048 3936
rect 278044 3952 278096 4004
rect 210792 3884 210844 3936
rect 219532 3884 219584 3936
rect 220728 3884 220780 3936
rect 225052 3884 225104 3936
rect 226248 3884 226300 3936
rect 241612 3884 241664 3936
rect 242808 3884 242860 3936
rect 247132 3884 247184 3936
rect 248328 3884 248380 3936
rect 258172 3884 258224 3936
rect 259368 3884 259420 3936
rect 274732 3884 274784 3936
rect 275928 3884 275980 3936
rect 280252 3884 280304 3936
rect 281448 3884 281500 3936
rect 291292 3952 291344 4004
rect 292488 3952 292540 4004
rect 295984 3952 296036 4004
rect 469128 3952 469180 4004
rect 490104 3884 490156 3936
rect 45192 3816 45244 3868
rect 58624 3816 58676 3868
rect 69480 3816 69532 3868
rect 86592 3816 86644 3868
rect 88340 3816 88392 3868
rect 99288 3816 99340 3868
rect 129004 3816 129056 3868
rect 164148 3816 164200 3868
rect 164332 3816 164384 3868
rect 165528 3816 165580 3868
rect 169024 3816 169076 3868
rect 412824 3816 412876 3868
rect 423772 3816 423824 3868
rect 424968 3816 425020 3868
rect 440332 3816 440384 3868
rect 441528 3816 441580 3868
rect 446404 3816 446456 3868
rect 35256 3748 35308 3800
rect 53104 3748 53156 3800
rect 66168 3748 66220 3800
rect 85764 3748 85816 3800
rect 92296 3748 92348 3800
rect 109224 3748 109276 3800
rect 119344 3748 119396 3800
rect 126888 3748 126940 3800
rect 127900 3748 127952 3800
rect 442632 3748 442684 3800
rect 445852 3748 445904 3800
rect 447048 3748 447100 3800
rect 523224 3748 523276 3800
rect 41880 3680 41932 3732
rect 83924 3680 83976 3732
rect 88616 3680 88668 3732
rect 102600 3680 102652 3732
rect 104440 3680 104492 3732
rect 123576 3680 123628 3732
rect 128084 3680 128136 3732
rect 456708 3680 456760 3732
rect 456892 3680 456944 3732
rect 458088 3680 458140 3732
rect 462412 3680 462464 3732
rect 463608 3680 463660 3732
rect 37464 3612 37516 3664
rect 83096 3612 83148 3664
rect 92112 3612 92164 3664
rect 125784 3612 125836 3664
rect 127992 3612 128044 3664
rect 476856 3680 476908 3732
rect 33048 3544 33100 3596
rect 75736 3544 75788 3596
rect 27528 3476 27580 3528
rect 31024 3476 31076 3528
rect 80060 3544 80112 3596
rect 29736 3408 29788 3460
rect 75920 3476 75972 3528
rect 77208 3476 77260 3528
rect 82728 3476 82780 3528
rect 87328 3544 87380 3596
rect 90732 3544 90784 3596
rect 86040 3476 86092 3528
rect 87236 3476 87288 3528
rect 89352 3476 89404 3528
rect 91560 3476 91612 3528
rect 91928 3544 91980 3596
rect 112536 3544 112588 3596
rect 121276 3544 121328 3596
rect 473544 3612 473596 3664
rect 473452 3544 473504 3596
rect 474648 3544 474700 3596
rect 484400 3544 484452 3596
rect 485688 3544 485740 3596
rect 115848 3476 115900 3528
rect 122564 3476 122616 3528
rect 493416 3544 493468 3596
rect 501052 3544 501104 3596
rect 502248 3544 502300 3596
rect 506572 3544 506624 3596
rect 507768 3544 507820 3596
rect 545212 3544 545264 3596
rect 546408 3544 546460 3596
rect 550732 3544 550784 3596
rect 551928 3544 551980 3596
rect 490012 3476 490064 3528
rect 491208 3476 491260 3528
rect 512000 3476 512052 3528
rect 513288 3476 513340 3528
rect 539600 3476 539652 3528
rect 540888 3476 540940 3528
rect 28632 3340 28684 3392
rect 83004 3408 83056 3460
rect 87420 3408 87472 3460
rect 90456 3408 90508 3460
rect 59360 3340 59412 3392
rect 60648 3340 60700 3392
rect 70400 3340 70452 3392
rect 71688 3340 71740 3392
rect 88524 3340 88576 3392
rect 92664 3340 92716 3392
rect 89812 3272 89864 3324
rect 118056 3408 118108 3460
rect 121552 3408 121604 3460
rect 496728 3408 496780 3460
rect 100024 3340 100076 3392
rect 101496 3340 101548 3392
rect 135904 3340 135956 3392
rect 137928 3340 137980 3392
rect 153200 3340 153252 3392
rect 154488 3340 154540 3392
rect 164148 3340 164200 3392
rect 167736 3340 167788 3392
rect 180800 3340 180852 3392
rect 182088 3340 182140 3392
rect 186320 3340 186372 3392
rect 187608 3340 187660 3392
rect 197360 3340 197412 3392
rect 198648 3340 198700 3392
rect 202880 3340 202932 3392
rect 204168 3340 204220 3392
rect 236000 3340 236052 3392
rect 237288 3340 237340 3392
rect 252560 3340 252612 3392
rect 253848 3340 253900 3392
rect 269120 3340 269172 3392
rect 270408 3340 270460 3392
rect 285680 3340 285732 3392
rect 286968 3340 287020 3392
rect 302240 3340 302292 3392
rect 303528 3340 303580 3392
rect 313280 3340 313332 3392
rect 314568 3340 314620 3392
rect 318800 3340 318852 3392
rect 320088 3340 320140 3392
rect 335360 3340 335412 3392
rect 336648 3340 336700 3392
rect 351920 3340 351972 3392
rect 353208 3340 353260 3392
rect 362960 3340 363012 3392
rect 364248 3340 364300 3392
rect 368480 3340 368532 3392
rect 369768 3340 369820 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 379520 3340 379572 3392
rect 380808 3340 380860 3392
rect 385040 3340 385092 3392
rect 386328 3340 386380 3392
rect 401600 3340 401652 3392
rect 402888 3340 402940 3392
rect 412732 3340 412784 3392
rect 413928 3340 413980 3392
rect 418160 3340 418212 3392
rect 419448 3340 419500 3392
rect 429200 3340 429252 3392
rect 430488 3340 430540 3392
rect 434720 3340 434772 3392
rect 436008 3340 436060 3392
rect 451280 3340 451332 3392
rect 452568 3340 452620 3392
rect 456708 3340 456760 3392
rect 459192 3340 459244 3392
rect 131764 3204 131816 3256
rect 133512 3204 133564 3256
rect 87144 3136 87196 3188
rect 89352 3136 89404 3188
rect 36360 3000 36412 3052
rect 43444 3000 43496 3052
rect 80520 2796 80572 2848
rect 82360 2796 82412 2848
rect 478880 1096 478932 1148
rect 480168 1096 480220 1148
rect 534080 688 534132 740
rect 535368 688 535420 740
<< metal2 >>
rect 9692 703582 10732 703610
rect 3422 694920 3478 694929
rect 3422 694855 3478 694864
rect 3436 694210 3464 694855
rect 3424 694204 3476 694210
rect 3424 694146 3476 694152
rect 3422 678192 3478 678201
rect 3422 678127 3478 678136
rect 3436 677618 3464 678127
rect 3424 677612 3476 677618
rect 3424 677554 3476 677560
rect 3422 661464 3478 661473
rect 3422 661399 3478 661408
rect 3436 661094 3464 661399
rect 3424 661088 3476 661094
rect 3424 661030 3476 661036
rect 3238 644736 3294 644745
rect 3238 644671 3294 644680
rect 3252 644502 3280 644671
rect 3240 644496 3292 644502
rect 3240 644438 3292 644444
rect 3422 628008 3478 628017
rect 3422 627943 3424 627952
rect 3476 627943 3478 627952
rect 3424 627914 3476 627920
rect 3422 611280 3478 611289
rect 3422 611215 3478 611224
rect 3436 610026 3464 611215
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3422 594552 3478 594561
rect 3422 594487 3478 594496
rect 3054 577824 3110 577833
rect 3054 577759 3110 577768
rect 3068 576910 3096 577759
rect 3056 576904 3108 576910
rect 3056 576846 3108 576852
rect 3054 561096 3110 561105
rect 3054 561031 3110 561040
rect 3068 560318 3096 561031
rect 3056 560312 3108 560318
rect 3056 560254 3108 560260
rect 3330 510912 3386 510921
rect 3330 510847 3386 510856
rect 3344 510678 3372 510847
rect 3332 510672 3384 510678
rect 3332 510614 3384 510620
rect 3330 494184 3386 494193
rect 3330 494119 3386 494128
rect 3344 494086 3372 494119
rect 3332 494080 3384 494086
rect 3332 494022 3384 494028
rect 3146 477456 3202 477465
rect 3146 477391 3202 477400
rect 3160 476202 3188 477391
rect 3148 476196 3200 476202
rect 3148 476138 3200 476144
rect 3146 460728 3202 460737
rect 3146 460663 3202 460672
rect 3160 459610 3188 460663
rect 3148 459604 3200 459610
rect 3148 459546 3200 459552
rect 3330 444000 3386 444009
rect 3330 443935 3386 443944
rect 3344 443018 3372 443935
rect 3332 443012 3384 443018
rect 3332 442954 3384 442960
rect 3330 427272 3386 427281
rect 3330 427207 3386 427216
rect 3344 426494 3372 427207
rect 3332 426488 3384 426494
rect 3332 426430 3384 426436
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3330 377088 3386 377097
rect 3330 377023 3386 377032
rect 3344 376786 3372 377023
rect 3332 376780 3384 376786
rect 3332 376722 3384 376728
rect 3330 360360 3386 360369
rect 3330 360295 3386 360304
rect 3344 360262 3372 360295
rect 3332 360256 3384 360262
rect 3332 360198 3384 360204
rect 3330 343632 3386 343641
rect 3330 343567 3386 343576
rect 3344 342310 3372 343567
rect 3332 342304 3384 342310
rect 3332 342246 3384 342252
rect 3330 326904 3386 326913
rect 3330 326839 3386 326848
rect 3344 325718 3372 326839
rect 3332 325712 3384 325718
rect 3332 325654 3384 325660
rect 3330 310176 3386 310185
rect 3330 310111 3386 310120
rect 3344 309194 3372 310111
rect 3332 309188 3384 309194
rect 3332 309130 3384 309136
rect 3330 293448 3386 293457
rect 3330 293383 3386 293392
rect 3344 292602 3372 293383
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3330 276720 3386 276729
rect 3330 276655 3386 276664
rect 3344 276078 3372 276655
rect 3332 276072 3384 276078
rect 3332 276014 3384 276020
rect 2962 259992 3018 260001
rect 2962 259927 3018 259936
rect 2976 259486 3004 259927
rect 2964 259480 3016 259486
rect 2964 259422 3016 259428
rect 3330 243264 3386 243273
rect 3330 243199 3386 243208
rect 3344 242962 3372 243199
rect 3332 242956 3384 242962
rect 3332 242898 3384 242904
rect 3330 226536 3386 226545
rect 3330 226471 3386 226480
rect 3344 226438 3372 226471
rect 3332 226432 3384 226438
rect 3332 226374 3384 226380
rect 3332 209840 3384 209846
rect 3330 209808 3332 209817
rect 3384 209808 3386 209817
rect 3330 209743 3386 209752
rect 3330 193080 3386 193089
rect 3330 193015 3386 193024
rect 3344 191894 3372 193015
rect 3332 191888 3384 191894
rect 3332 191830 3384 191836
rect 3054 176352 3110 176361
rect 3054 176287 3110 176296
rect 3068 175302 3096 176287
rect 3056 175296 3108 175302
rect 3056 175238 3108 175244
rect 3146 159624 3202 159633
rect 3146 159559 3202 159568
rect 3160 158778 3188 159559
rect 3148 158772 3200 158778
rect 3148 158714 3200 158720
rect 3436 155582 3464 594487
rect 3514 544368 3570 544377
rect 3514 544303 3570 544312
rect 3424 155576 3476 155582
rect 3424 155518 3476 155524
rect 3528 155514 3556 544303
rect 3606 527640 3662 527649
rect 3606 527575 3662 527584
rect 3620 527202 3648 527575
rect 3608 527196 3660 527202
rect 3608 527138 3660 527144
rect 3606 393816 3662 393825
rect 3606 393751 3662 393760
rect 3620 393378 3648 393751
rect 3608 393372 3660 393378
rect 3608 393314 3660 393320
rect 9692 156874 9720 703582
rect 10704 703474 10732 703582
rect 10846 703520 10958 704960
rect 32466 703520 32578 704960
rect 54086 703520 54198 704960
rect 75706 703520 75818 704960
rect 97326 703520 97438 704960
rect 118946 703520 119058 704960
rect 139412 703582 140452 703610
rect 10888 703474 10916 703520
rect 10704 703446 10916 703474
rect 32508 700670 32536 703520
rect 54128 702434 54156 703520
rect 75748 703050 75776 703520
rect 74540 703044 74592 703050
rect 74540 702986 74592 702992
rect 75736 703044 75788 703050
rect 75736 702986 75788 702992
rect 53852 702406 54156 702434
rect 32496 700664 32548 700670
rect 32496 700606 32548 700612
rect 9680 156868 9732 156874
rect 9680 156810 9732 156816
rect 3516 155508 3568 155514
rect 3516 155450 3568 155456
rect 53852 154222 53880 702406
rect 74552 157010 74580 702986
rect 97368 700806 97396 703520
rect 118988 702434 119016 703520
rect 118712 702406 119016 702434
rect 97356 700800 97408 700806
rect 97356 700742 97408 700748
rect 109040 700800 109092 700806
rect 109040 700742 109092 700748
rect 107660 700732 107712 700738
rect 107660 700674 107712 700680
rect 106280 700528 106332 700534
rect 106280 700470 106332 700476
rect 103520 700460 103572 700466
rect 103520 700402 103572 700408
rect 102140 700392 102192 700398
rect 102140 700334 102192 700340
rect 100852 695564 100904 695570
rect 100852 695506 100904 695512
rect 100208 663808 100260 663814
rect 100208 663750 100260 663756
rect 99656 648644 99708 648650
rect 99656 648586 99708 648592
rect 99472 616888 99524 616894
rect 99472 616830 99524 616836
rect 98552 601724 98604 601730
rect 98552 601666 98604 601672
rect 98276 586560 98328 586566
rect 98276 586502 98328 586508
rect 97448 554804 97500 554810
rect 97448 554746 97500 554752
rect 96896 539640 96948 539646
rect 96896 539582 96948 539588
rect 95792 507884 95844 507890
rect 95792 507826 95844 507832
rect 95516 476128 95568 476134
rect 95516 476070 95568 476076
rect 95332 460964 95384 460970
rect 95332 460906 95384 460912
rect 94688 429208 94740 429214
rect 94688 429150 94740 429156
rect 94136 414044 94188 414050
rect 94136 413986 94188 413992
rect 93952 382288 94004 382294
rect 93952 382230 94004 382236
rect 92480 367124 92532 367130
rect 92480 367066 92532 367072
rect 91100 320204 91152 320210
rect 91100 320146 91152 320152
rect 89720 273284 89772 273290
rect 89720 273226 89772 273232
rect 88340 194608 88392 194614
rect 88340 194550 88392 194556
rect 88352 160274 88380 194550
rect 88616 179444 88668 179450
rect 88616 179386 88668 179392
rect 88340 160268 88392 160274
rect 88340 160210 88392 160216
rect 74540 157004 74592 157010
rect 74540 156946 74592 156952
rect 53840 154216 53892 154222
rect 53840 154158 53892 154164
rect 7564 152720 7616 152726
rect 7564 152662 7616 152668
rect 4804 152448 4856 152454
rect 4804 152390 4856 152396
rect 3792 152380 3844 152386
rect 3792 152322 3844 152328
rect 3516 151156 3568 151162
rect 3516 151098 3568 151104
rect 3240 150544 3292 150550
rect 3240 150486 3292 150492
rect 3252 142202 3280 150486
rect 3424 149388 3476 149394
rect 3424 149330 3476 149336
rect 3436 142905 3464 149330
rect 3422 142896 3478 142905
rect 3422 142831 3478 142840
rect 3252 142174 3464 142202
rect 3332 126472 3384 126478
rect 3332 126414 3384 126420
rect 3344 126177 3372 126414
rect 3330 126168 3386 126177
rect 3330 126103 3386 126112
rect 2780 110152 2832 110158
rect 2780 110094 2832 110100
rect 2792 109449 2820 110094
rect 2778 109440 2834 109449
rect 2778 109375 2834 109384
rect 3436 9081 3464 142174
rect 3528 25809 3556 151098
rect 3700 150680 3752 150686
rect 3700 150622 3752 150628
rect 3608 150612 3660 150618
rect 3608 150554 3660 150560
rect 3620 42537 3648 150554
rect 3712 59265 3740 150622
rect 3804 75993 3832 152322
rect 3884 150748 3936 150754
rect 3884 150690 3936 150696
rect 3896 92721 3924 150690
rect 4816 110158 4844 152390
rect 7576 126478 7604 152662
rect 81900 152584 81952 152590
rect 81900 152526 81952 152532
rect 86866 152552 86922 152561
rect 80888 152516 80940 152522
rect 80888 152458 80940 152464
rect 7564 126472 7616 126478
rect 7564 126414 7616 126420
rect 4804 110152 4856 110158
rect 4804 110094 4856 110100
rect 80900 100230 80928 152458
rect 81716 152176 81768 152182
rect 81716 152118 81768 152124
rect 81440 152108 81492 152114
rect 81440 152050 81492 152056
rect 80980 150204 81032 150210
rect 80980 150146 81032 150152
rect 80888 100224 80940 100230
rect 80888 100166 80940 100172
rect 77852 100088 77904 100094
rect 77852 100030 77904 100036
rect 64880 97708 64932 97714
rect 64880 97650 64932 97656
rect 62764 97640 62816 97646
rect 62764 97582 62816 97588
rect 58624 97572 58676 97578
rect 58624 97514 58676 97520
rect 53104 97504 53156 97510
rect 53104 97446 53156 97452
rect 43444 97368 43496 97374
rect 43444 97310 43496 97316
rect 31024 97300 31076 97306
rect 31024 97242 31076 97248
rect 3882 92712 3938 92721
rect 3882 92647 3938 92656
rect 3790 75984 3846 75993
rect 3790 75919 3846 75928
rect 3698 59256 3754 59265
rect 3698 59191 3754 59200
rect 30380 44872 30432 44878
rect 30380 44814 30432 44820
rect 3606 42528 3662 42537
rect 3606 42463 3662 42472
rect 3514 25800 3570 25809
rect 3514 25735 3570 25744
rect 30392 16574 30420 44814
rect 30392 16546 30880 16574
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 26424 7608 26476 7614
rect 26424 7550 26476 7556
rect 25320 4956 25372 4962
rect 25320 4898 25372 4904
rect 24216 4888 24268 4894
rect 24216 4830 24268 4836
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23124 480 23152 4762
rect 24228 480 24256 4830
rect 25332 480 25360 4898
rect 26436 480 26464 7550
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27540 480 27568 3470
rect 29736 3460 29788 3466
rect 29736 3402 29788 3408
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28644 480 28672 3334
rect 29748 480 29776 3402
rect 30852 480 30880 16546
rect 31036 3534 31064 97242
rect 40040 87644 40092 87650
rect 40040 87586 40092 87592
rect 31760 84924 31812 84930
rect 31760 84866 31812 84872
rect 31772 16574 31800 84866
rect 38660 21412 38712 21418
rect 38660 21354 38712 21360
rect 38672 16574 38700 21354
rect 40052 16574 40080 87586
rect 31772 16546 31984 16574
rect 38672 16546 39712 16574
rect 40052 16546 40816 16574
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31956 480 31984 16546
rect 38568 6248 38620 6254
rect 38568 6190 38620 6196
rect 34152 6180 34204 6186
rect 34152 6122 34204 6128
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33060 480 33088 3538
rect 34164 480 34192 6122
rect 35256 3800 35308 3806
rect 35256 3742 35308 3748
rect 35268 480 35296 3742
rect 37464 3664 37516 3670
rect 37464 3606 37516 3612
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36372 480 36400 2994
rect 37476 480 37504 3606
rect 38580 480 38608 6190
rect 39684 480 39712 16546
rect 40788 480 40816 16546
rect 42982 7576 43038 7585
rect 42982 7511 43038 7520
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41892 480 41920 3674
rect 42996 480 43024 7511
rect 43456 3058 43484 97310
rect 46940 44940 46992 44946
rect 46940 44882 46992 44888
rect 46952 16574 46980 44882
rect 46952 16546 47440 16574
rect 46294 4856 46350 4865
rect 46294 4791 46350 4800
rect 44088 3936 44140 3942
rect 44088 3878 44140 3884
rect 43444 3052 43496 3058
rect 43444 2994 43496 3000
rect 44100 480 44128 3878
rect 45192 3868 45244 3874
rect 45192 3810 45244 3816
rect 45204 480 45232 3810
rect 46308 480 46336 4791
rect 47412 480 47440 16546
rect 48504 6316 48556 6322
rect 48504 6258 48556 6264
rect 48516 480 48544 6258
rect 52920 5160 52972 5166
rect 52920 5102 52972 5108
rect 50712 5092 50764 5098
rect 50712 5034 50764 5040
rect 49608 5024 49660 5030
rect 49608 4966 49660 4972
rect 49620 480 49648 4966
rect 50724 480 50752 5034
rect 51816 4004 51868 4010
rect 51816 3946 51868 3952
rect 51828 480 51856 3946
rect 52932 480 52960 5102
rect 53116 3806 53144 97446
rect 54484 97436 54536 97442
rect 54484 97378 54536 97384
rect 53840 86284 53892 86290
rect 53840 86226 53892 86232
rect 53852 16574 53880 86226
rect 53852 16546 54064 16574
rect 53104 3800 53156 3806
rect 53104 3742 53156 3748
rect 54036 480 54064 16546
rect 54496 3942 54524 97378
rect 56600 87712 56652 87718
rect 56600 87654 56652 87660
rect 56612 16574 56640 87654
rect 56612 16546 57376 16574
rect 55128 6384 55180 6390
rect 55128 6326 55180 6332
rect 54484 3936 54536 3942
rect 54484 3878 54536 3884
rect 55140 480 55168 6326
rect 56232 5228 56284 5234
rect 56232 5170 56284 5176
rect 56244 480 56272 5170
rect 57348 480 57376 16546
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 58452 480 58480 3878
rect 58636 3874 58664 97514
rect 59358 87544 59414 87553
rect 59358 87479 59414 87488
rect 58624 3868 58676 3874
rect 58624 3810 58676 3816
rect 59372 3398 59400 87479
rect 61752 7676 61804 7682
rect 61752 7618 61804 7624
rect 59542 4992 59598 5001
rect 59542 4927 59598 4936
rect 59360 3392 59412 3398
rect 59360 3334 59412 3340
rect 59556 480 59584 4927
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60660 480 60688 3334
rect 61764 480 61792 7618
rect 62776 4010 62804 97582
rect 64892 16574 64920 97650
rect 77864 97442 77892 100030
rect 80428 100020 80480 100026
rect 80428 99962 80480 99968
rect 79784 99748 79836 99754
rect 79784 99690 79836 99696
rect 79796 97510 79824 99690
rect 79784 97504 79836 97510
rect 79784 97446 79836 97452
rect 77852 97436 77904 97442
rect 77852 97378 77904 97384
rect 80440 97374 80468 99962
rect 80428 97368 80480 97374
rect 80428 97310 80480 97316
rect 71044 97028 71096 97034
rect 71044 96970 71096 96976
rect 70400 45008 70452 45014
rect 70400 44950 70452 44956
rect 64892 16546 65104 16574
rect 63960 6520 64012 6526
rect 63960 6462 64012 6468
rect 62856 6452 62908 6458
rect 62856 6394 62908 6400
rect 62764 4004 62816 4010
rect 62764 3946 62816 3952
rect 62868 480 62896 6394
rect 63972 480 64000 6462
rect 65076 480 65104 16546
rect 68376 6656 68428 6662
rect 68376 6598 68428 6604
rect 67272 6588 67324 6594
rect 67272 6530 67324 6536
rect 66168 3800 66220 3806
rect 66168 3742 66220 3748
rect 66180 480 66208 3742
rect 67284 480 67312 6530
rect 68388 480 68416 6598
rect 69480 3868 69532 3874
rect 69480 3810 69532 3816
rect 69492 480 69520 3810
rect 70412 3398 70440 44950
rect 70584 6724 70636 6730
rect 70584 6666 70636 6672
rect 70400 3392 70452 3398
rect 70400 3334 70452 3340
rect 70596 480 70624 6666
rect 71056 3942 71084 96970
rect 80992 96354 81020 150146
rect 81348 150000 81400 150006
rect 81348 149942 81400 149948
rect 81164 149932 81216 149938
rect 81164 149874 81216 149880
rect 81072 149796 81124 149802
rect 81072 149738 81124 149744
rect 80980 96348 81032 96354
rect 80980 96290 81032 96296
rect 81084 95810 81112 149738
rect 81176 95878 81204 149874
rect 81256 149728 81308 149734
rect 81256 149670 81308 149676
rect 81268 96082 81296 149670
rect 81360 96422 81388 149942
rect 81452 113174 81480 152050
rect 81452 113146 81572 113174
rect 81544 109034 81572 113146
rect 81452 109006 81572 109034
rect 81728 109018 81756 152118
rect 81808 149592 81860 149598
rect 81808 149534 81860 149540
rect 81452 99958 81480 109006
rect 81636 108990 81756 109018
rect 81636 106274 81664 108990
rect 81636 106246 81756 106274
rect 81530 104408 81586 104417
rect 81530 104343 81586 104352
rect 81440 99952 81492 99958
rect 81440 99894 81492 99900
rect 81440 99816 81492 99822
rect 81440 99758 81492 99764
rect 81348 96416 81400 96422
rect 81348 96358 81400 96364
rect 81452 96286 81480 99758
rect 81544 97238 81572 104343
rect 81624 99884 81676 99890
rect 81624 99826 81676 99832
rect 81532 97232 81584 97238
rect 81532 97174 81584 97180
rect 81440 96280 81492 96286
rect 81440 96222 81492 96228
rect 81256 96076 81308 96082
rect 81256 96018 81308 96024
rect 81164 95872 81216 95878
rect 81164 95814 81216 95820
rect 81072 95804 81124 95810
rect 81072 95746 81124 95752
rect 81532 94716 81584 94722
rect 81532 94658 81584 94664
rect 77300 87780 77352 87786
rect 77300 87722 77352 87728
rect 75920 83496 75972 83502
rect 75920 83438 75972 83444
rect 73896 6792 73948 6798
rect 73896 6734 73948 6740
rect 71044 3936 71096 3942
rect 71044 3878 71096 3884
rect 72792 3936 72844 3942
rect 72792 3878 72844 3884
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71700 480 71728 3334
rect 72804 480 72832 3878
rect 73908 480 73936 6734
rect 75000 5364 75052 5370
rect 75000 5306 75052 5312
rect 75012 480 75040 5306
rect 75736 4140 75788 4146
rect 75736 4082 75788 4088
rect 75748 3602 75776 4082
rect 75736 3596 75788 3602
rect 75736 3538 75788 3544
rect 75932 3534 75960 83438
rect 77312 16574 77340 87722
rect 77312 16546 78352 16574
rect 76104 4004 76156 4010
rect 76104 3946 76156 3952
rect 75920 3528 75972 3534
rect 75920 3470 75972 3476
rect 76116 480 76144 3946
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 77220 480 77248 3470
rect 78324 480 78352 16546
rect 80060 5296 80112 5302
rect 80060 5238 80112 5244
rect 79416 4072 79468 4078
rect 79416 4014 79468 4020
rect 79428 480 79456 4014
rect 80072 3602 80100 5238
rect 81544 4826 81572 94658
rect 81636 4894 81664 99826
rect 81728 99278 81756 106246
rect 81820 104417 81848 149534
rect 81806 104408 81862 104417
rect 81806 104343 81862 104352
rect 81912 104258 81940 152526
rect 86866 152487 86922 152496
rect 82360 152312 82412 152318
rect 82360 152254 82412 152260
rect 82176 152244 82228 152250
rect 82176 152186 82228 152192
rect 81992 149524 82044 149530
rect 81992 149466 82044 149472
rect 81820 104230 81940 104258
rect 81820 100298 81848 104230
rect 81900 101516 81952 101522
rect 81900 101458 81952 101464
rect 81808 100292 81860 100298
rect 81808 100234 81860 100240
rect 81808 100156 81860 100162
rect 81808 100098 81860 100104
rect 81716 99272 81768 99278
rect 81716 99214 81768 99220
rect 81820 97714 81848 100098
rect 81912 99822 81940 101458
rect 81900 99816 81952 99822
rect 81900 99758 81952 99764
rect 82004 97782 82032 149466
rect 82084 149456 82136 149462
rect 82084 149398 82136 149404
rect 82096 97850 82124 149398
rect 82084 97844 82136 97850
rect 82084 97786 82136 97792
rect 81992 97776 82044 97782
rect 81992 97718 82044 97724
rect 81808 97708 81860 97714
rect 81808 97650 81860 97656
rect 81808 97096 81860 97102
rect 81808 97038 81860 97044
rect 81624 4888 81676 4894
rect 81624 4830 81676 4836
rect 81532 4820 81584 4826
rect 81532 4762 81584 4768
rect 80060 3596 80112 3602
rect 80060 3538 80112 3544
rect 80520 2848 80572 2854
rect 80520 2790 80572 2796
rect 80532 480 80560 2790
rect 21978 -960 22090 480
rect 23082 -960 23194 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26394 -960 26506 480
rect 27498 -960 27610 480
rect 28602 -960 28714 480
rect 29706 -960 29818 480
rect 30810 -960 30922 480
rect 31914 -960 32026 480
rect 33018 -960 33130 480
rect 34122 -960 34234 480
rect 35226 -960 35338 480
rect 36330 -960 36442 480
rect 37434 -960 37546 480
rect 38538 -960 38650 480
rect 39642 -960 39754 480
rect 40746 -960 40858 480
rect 41850 -960 41962 480
rect 42954 -960 43066 480
rect 44058 -960 44170 480
rect 45162 -960 45274 480
rect 46266 -960 46378 480
rect 47370 -960 47482 480
rect 48474 -960 48586 480
rect 49578 -960 49690 480
rect 50682 -960 50794 480
rect 51786 -960 51898 480
rect 52890 -960 53002 480
rect 53994 -960 54106 480
rect 55098 -960 55210 480
rect 56202 -960 56314 480
rect 57306 -960 57418 480
rect 58410 -960 58522 480
rect 59514 -960 59626 480
rect 60618 -960 60730 480
rect 61722 -960 61834 480
rect 62826 -960 62938 480
rect 63930 -960 64042 480
rect 65034 -960 65146 480
rect 66138 -960 66250 480
rect 67242 -960 67354 480
rect 68346 -960 68458 480
rect 69450 -960 69562 480
rect 70554 -960 70666 480
rect 71658 -960 71770 480
rect 72762 -960 72874 480
rect 73866 -960 73978 480
rect 74970 -960 75082 480
rect 76074 -960 76186 480
rect 77178 -960 77290 480
rect 78282 -960 78394 480
rect 79386 -960 79498 480
rect 80490 -960 80602 480
rect 81594 354 81706 480
rect 81820 354 81848 97038
rect 82188 96966 82216 152186
rect 82268 151836 82320 151842
rect 82268 151778 82320 151784
rect 82176 96960 82228 96966
rect 82176 96902 82228 96908
rect 82280 96558 82308 151778
rect 82372 101522 82400 152254
rect 85856 152040 85908 152046
rect 85856 151982 85908 151988
rect 85486 150512 85542 150521
rect 85486 150447 85542 150456
rect 85500 149954 85528 150447
rect 85868 149954 85896 151982
rect 86880 149954 86908 152487
rect 88062 152416 88118 152425
rect 88062 152351 88118 152360
rect 87788 150816 87840 150822
rect 87788 150758 87840 150764
rect 87800 149954 87828 150758
rect 88076 149954 88104 152351
rect 88524 150476 88576 150482
rect 88524 150418 88576 150424
rect 88536 149954 88564 150418
rect 85468 149926 85528 149954
rect 85744 149926 85896 149954
rect 86848 149926 86908 149954
rect 87676 149926 87828 149954
rect 87952 149926 88104 149954
rect 88504 149926 88564 149954
rect 88628 149954 88656 179386
rect 88892 164280 88944 164286
rect 88892 164222 88944 164228
rect 88904 149954 88932 164222
rect 89444 160268 89496 160274
rect 89444 160210 89496 160216
rect 89456 149954 89484 160210
rect 89732 153270 89760 273226
rect 89996 241528 90048 241534
rect 89996 241470 90048 241476
rect 89812 226364 89864 226370
rect 89812 226306 89864 226312
rect 89720 153264 89772 153270
rect 89720 153206 89772 153212
rect 89824 150226 89852 226306
rect 90008 153338 90036 241470
rect 90088 211200 90140 211206
rect 90088 211142 90140 211148
rect 89996 153332 90048 153338
rect 89996 153274 90048 153280
rect 90100 150226 90128 211142
rect 90548 153332 90600 153338
rect 90548 153274 90600 153280
rect 89824 150198 89898 150226
rect 90100 150198 90174 150226
rect 88628 149926 88780 149954
rect 88904 149926 89056 149954
rect 89456 149926 89608 149954
rect 89870 149940 89898 150198
rect 90146 149940 90174 150198
rect 90560 149954 90588 153274
rect 91112 153270 91140 320146
rect 91376 305040 91428 305046
rect 91376 304982 91428 304988
rect 91192 258120 91244 258126
rect 91192 258062 91244 258068
rect 90824 153264 90876 153270
rect 90824 153206 90876 153212
rect 91100 153264 91152 153270
rect 91100 153206 91152 153212
rect 90836 149954 90864 153206
rect 91204 150226 91232 258062
rect 91388 153338 91416 304982
rect 91652 288448 91704 288454
rect 91652 288390 91704 288396
rect 91376 153332 91428 153338
rect 91376 153274 91428 153280
rect 91204 150198 91278 150226
rect 90560 149926 90712 149954
rect 90836 149926 90988 149954
rect 91250 149940 91278 150198
rect 91514 150204 91566 150210
rect 91514 150146 91566 150152
rect 91526 149940 91554 150146
rect 91664 149954 91692 288390
rect 92492 153338 92520 367066
rect 92756 351960 92808 351966
rect 92756 351902 92808 351908
rect 92768 159254 92796 351902
rect 92848 335368 92900 335374
rect 92848 335310 92900 335316
rect 92756 159248 92808 159254
rect 92756 159190 92808 159196
rect 92204 153332 92256 153338
rect 92204 153274 92256 153280
rect 92480 153332 92532 153338
rect 92480 153274 92532 153280
rect 91928 153264 91980 153270
rect 91928 153206 91980 153212
rect 91940 149954 91968 153206
rect 92216 149954 92244 153274
rect 92860 150226 92888 335310
rect 93308 159248 93360 159254
rect 93308 159190 93360 159196
rect 93032 153332 93084 153338
rect 93032 153274 93084 153280
rect 92860 150198 92934 150226
rect 91664 149926 91816 149954
rect 91940 149926 92092 149954
rect 92216 149926 92368 149954
rect 92906 149940 92934 150198
rect 93044 149954 93072 153274
rect 93320 149954 93348 159190
rect 93964 150226 93992 382230
rect 93964 150198 94038 150226
rect 93044 149926 93196 149954
rect 93320 149926 93472 149954
rect 94010 149940 94038 150198
rect 94148 149954 94176 413986
rect 94412 398880 94464 398886
rect 94412 398822 94464 398828
rect 94424 149954 94452 398822
rect 94700 171134 94728 429150
rect 94700 171106 95004 171134
rect 94688 152516 94740 152522
rect 94688 152458 94740 152464
rect 94700 149954 94728 152458
rect 94976 149954 95004 171106
rect 95240 152040 95292 152046
rect 95240 151982 95292 151988
rect 95252 151094 95280 151982
rect 95240 151088 95292 151094
rect 95240 151030 95292 151036
rect 95344 150226 95372 460906
rect 95528 153338 95556 476070
rect 95608 445800 95660 445806
rect 95608 445742 95660 445748
rect 95516 153332 95568 153338
rect 95516 153274 95568 153280
rect 95620 150226 95648 445742
rect 95804 171134 95832 507826
rect 96712 492720 96764 492726
rect 96712 492662 96764 492668
rect 95804 171106 96384 171134
rect 96068 153332 96120 153338
rect 96068 153274 96120 153280
rect 95792 152584 95844 152590
rect 95792 152526 95844 152532
rect 95344 150198 95418 150226
rect 95620 150198 95694 150226
rect 94148 149926 94300 149954
rect 94424 149926 94576 149954
rect 94700 149926 94852 149954
rect 94976 149926 95128 149954
rect 95390 149940 95418 150198
rect 95666 149940 95694 150198
rect 95804 149954 95832 152526
rect 96080 149954 96108 153274
rect 96356 149954 96384 171106
rect 96724 150226 96752 492662
rect 96908 153338 96936 539582
rect 97172 523048 97224 523054
rect 97172 522990 97224 522996
rect 96896 153332 96948 153338
rect 96896 153274 96948 153280
rect 96896 152244 96948 152250
rect 96896 152186 96948 152192
rect 96724 150198 96798 150226
rect 95804 149926 95956 149954
rect 96080 149926 96232 149954
rect 96356 149926 96508 149954
rect 96770 149940 96798 150198
rect 96908 149954 96936 152186
rect 97184 149954 97212 522990
rect 97460 149954 97488 554746
rect 98288 153338 98316 586502
rect 98368 569968 98420 569974
rect 98368 569910 98420 569916
rect 97724 153332 97776 153338
rect 97724 153274 97776 153280
rect 98276 153332 98328 153338
rect 98276 153274 98328 153280
rect 97736 149954 97764 153274
rect 97998 152144 98054 152153
rect 97998 152079 98054 152088
rect 98012 151162 98040 152079
rect 98184 151836 98236 151842
rect 98184 151778 98236 151784
rect 98000 151156 98052 151162
rect 98000 151098 98052 151104
rect 98196 149954 98224 151778
rect 98380 150226 98408 569910
rect 98380 150198 98454 150226
rect 96908 149926 97060 149954
rect 97184 149926 97336 149954
rect 97460 149926 97612 149954
rect 97736 149926 97888 149954
rect 98164 149926 98224 149954
rect 98426 149940 98454 150198
rect 98564 149954 98592 601666
rect 98828 153332 98880 153338
rect 98828 153274 98880 153280
rect 98840 149954 98868 153274
rect 99104 152176 99156 152182
rect 99104 152118 99156 152124
rect 99116 149954 99144 152118
rect 99484 150226 99512 616830
rect 99484 150198 99558 150226
rect 98564 149926 98716 149954
rect 98840 149926 98992 149954
rect 99116 149926 99268 149954
rect 99530 149940 99558 150198
rect 99668 149954 99696 648586
rect 99932 633480 99984 633486
rect 99932 633422 99984 633428
rect 99944 149954 99972 633422
rect 100220 171134 100248 663750
rect 100220 171106 100524 171134
rect 100208 152108 100260 152114
rect 100208 152050 100260 152056
rect 100220 149954 100248 152050
rect 100496 149954 100524 171106
rect 100864 150226 100892 695506
rect 101036 680400 101088 680406
rect 101036 680342 101088 680348
rect 100864 150198 100938 150226
rect 99668 149926 99820 149954
rect 99944 149926 100096 149954
rect 100220 149926 100372 149954
rect 100496 149926 100648 149954
rect 100910 149940 100938 150198
rect 101048 149954 101076 680342
rect 102152 158302 102180 700334
rect 102232 700324 102284 700330
rect 102232 700266 102284 700272
rect 102140 158296 102192 158302
rect 102140 158238 102192 158244
rect 101864 155236 101916 155242
rect 101864 155178 101916 155184
rect 101772 153876 101824 153882
rect 101772 153818 101824 153824
rect 101312 152312 101364 152318
rect 101312 152254 101364 152260
rect 101324 149954 101352 152254
rect 101784 149954 101812 153818
rect 101048 149926 101200 149954
rect 101324 149926 101476 149954
rect 101752 149926 101812 149954
rect 101876 149954 101904 155178
rect 102244 150226 102272 700266
rect 103532 171134 103560 700402
rect 106292 171134 106320 700470
rect 103532 171106 104388 171134
rect 106292 171106 106596 171134
rect 103244 158296 103296 158302
rect 103244 158238 103296 158244
rect 102968 155304 103020 155310
rect 102968 155246 103020 155252
rect 102876 153944 102928 153950
rect 102876 153886 102928 153892
rect 102690 152280 102746 152289
rect 102690 152215 102746 152224
rect 102244 150198 102318 150226
rect 101876 149926 102028 149954
rect 102290 149940 102318 150198
rect 102704 149954 102732 152215
rect 102888 149954 102916 153886
rect 102580 149926 102732 149954
rect 102856 149926 102916 149954
rect 102980 149954 103008 155246
rect 103256 149954 103284 158238
rect 104072 155372 104124 155378
rect 104072 155314 104124 155320
rect 103980 154012 104032 154018
rect 103980 153954 104032 153960
rect 103796 152040 103848 152046
rect 103796 151982 103848 151988
rect 103808 149954 103836 151982
rect 103992 149954 104020 153954
rect 102980 149926 103132 149954
rect 103256 149926 103408 149954
rect 103684 149926 103836 149954
rect 103960 149926 104020 149954
rect 104084 149954 104112 155314
rect 104360 149954 104388 171106
rect 106372 156800 106424 156806
rect 106372 156742 106424 156748
rect 105084 156732 105136 156738
rect 105084 156674 105136 156680
rect 104992 154080 105044 154086
rect 104992 154022 105044 154028
rect 104808 152108 104860 152114
rect 104808 152050 104860 152056
rect 104820 149954 104848 152050
rect 105004 150226 105032 154022
rect 105096 151814 105124 156674
rect 105452 156664 105504 156670
rect 105452 156606 105504 156612
rect 105096 151786 105216 151814
rect 105004 150198 105078 150226
rect 104084 149926 104236 149954
rect 104360 149926 104512 149954
rect 104788 149926 104848 149954
rect 105050 149940 105078 150198
rect 105188 149954 105216 151786
rect 105464 149954 105492 156606
rect 106188 154148 106240 154154
rect 106188 154090 106240 154096
rect 105726 151872 105782 151881
rect 105726 151807 105782 151816
rect 105740 149954 105768 151807
rect 106200 149954 106228 154090
rect 106384 150226 106412 156742
rect 106384 150198 106458 150226
rect 105188 149926 105340 149954
rect 105464 149926 105616 149954
rect 105740 149926 105892 149954
rect 106168 149926 106228 149954
rect 106430 149940 106458 150198
rect 106568 149954 106596 171106
rect 107672 158914 107700 700674
rect 107752 700596 107804 700602
rect 107752 700538 107804 700544
rect 107660 158908 107712 158914
rect 107660 158850 107712 158856
rect 107384 156936 107436 156942
rect 107384 156878 107436 156884
rect 107108 155440 107160 155446
rect 107108 155382 107160 155388
rect 106830 152008 106886 152017
rect 106830 151943 106886 151952
rect 106844 149954 106872 151943
rect 107120 149954 107148 155382
rect 107396 149954 107424 156878
rect 107764 150226 107792 700538
rect 109052 171134 109080 700742
rect 110972 700664 111024 700670
rect 110972 700606 111024 700612
rect 109052 171106 109908 171134
rect 108764 158908 108816 158914
rect 108764 158850 108816 158856
rect 108488 157072 108540 157078
rect 108488 157014 108540 157020
rect 108212 155644 108264 155650
rect 108212 155586 108264 155592
rect 108120 152244 108172 152250
rect 108120 152186 108172 152192
rect 107764 150198 107838 150226
rect 106568 149926 106720 149954
rect 106844 149926 106996 149954
rect 107120 149926 107272 149954
rect 107396 149926 107548 149954
rect 107810 149940 107838 150198
rect 108132 149954 108160 152186
rect 108100 149926 108160 149954
rect 108224 149954 108252 155586
rect 108500 149954 108528 157014
rect 108776 149954 108804 158850
rect 109684 157004 109736 157010
rect 109684 156946 109736 156952
rect 109592 154284 109644 154290
rect 109592 154226 109644 154232
rect 109316 152924 109368 152930
rect 109316 152866 109368 152872
rect 109328 149954 109356 152866
rect 109604 149954 109632 154226
rect 109696 150226 109724 156946
rect 109696 150198 109770 150226
rect 108224 149926 108376 149954
rect 108500 149926 108652 149954
rect 108776 149926 108928 149954
rect 109204 149926 109356 149954
rect 109480 149926 109632 149954
rect 109742 149940 109770 150198
rect 109880 149954 109908 171106
rect 110696 156868 110748 156874
rect 110696 156810 110748 156816
rect 110420 154216 110472 154222
rect 110420 154158 110472 154164
rect 110326 152688 110382 152697
rect 110326 152623 110382 152632
rect 110340 149954 110368 152623
rect 109880 149926 110032 149954
rect 110308 149926 110368 149954
rect 110432 149954 110460 154158
rect 110708 149954 110736 156810
rect 110984 149954 111012 700606
rect 111248 694204 111300 694210
rect 111248 694146 111300 694152
rect 111064 610020 111116 610026
rect 111064 609962 111116 609968
rect 111076 153202 111104 609962
rect 111260 171134 111288 694146
rect 112168 677612 112220 677618
rect 112168 677554 112220 677560
rect 111892 661088 111944 661094
rect 111892 661030 111944 661036
rect 111260 171106 111564 171134
rect 111064 153196 111116 153202
rect 111064 153138 111116 153144
rect 111432 152176 111484 152182
rect 111432 152118 111484 152124
rect 111444 149954 111472 152118
rect 110432 149926 110584 149954
rect 110708 149926 110860 149954
rect 110984 149926 111136 149954
rect 111412 149926 111472 149954
rect 111536 149954 111564 171106
rect 111904 150226 111932 661030
rect 112180 150226 112208 677554
rect 112352 644496 112404 644502
rect 112352 644438 112404 644444
rect 111904 150198 111978 150226
rect 112180 150198 112254 150226
rect 111536 149926 111688 149954
rect 111950 149940 111978 150198
rect 112226 149940 112254 150198
rect 112364 149870 112392 644438
rect 113364 627972 113416 627978
rect 113364 627914 113416 627920
rect 112444 560312 112496 560318
rect 112444 560254 112496 560260
rect 112456 151910 112484 560254
rect 112536 510672 112588 510678
rect 112536 510614 112588 510620
rect 112444 151904 112496 151910
rect 112444 151846 112496 151852
rect 112548 151842 112576 510614
rect 112904 153196 112956 153202
rect 112904 153138 112956 153144
rect 112626 152008 112682 152017
rect 112626 151943 112682 151952
rect 112536 151836 112588 151842
rect 112536 151778 112588 151784
rect 112640 149954 112668 151943
rect 112516 149926 112668 149954
rect 112916 149954 112944 153138
rect 113376 149954 113404 627914
rect 114008 576904 114060 576910
rect 114008 576846 114060 576852
rect 113824 459604 113876 459610
rect 113824 459546 113876 459552
rect 113732 155576 113784 155582
rect 113732 155518 113784 155524
rect 113640 151972 113692 151978
rect 113640 151914 113692 151920
rect 113652 149954 113680 151914
rect 112916 149926 113068 149954
rect 113344 149926 113404 149954
rect 113620 149926 113680 149954
rect 113744 149954 113772 155518
rect 113836 153202 113864 459546
rect 113916 409896 113968 409902
rect 113916 409838 113968 409844
rect 113928 155922 113956 409838
rect 114020 171134 114048 576846
rect 115112 527196 115164 527202
rect 115112 527138 115164 527144
rect 114020 171106 114324 171134
rect 113916 155916 113968 155922
rect 113916 155858 113968 155864
rect 113824 153196 113876 153202
rect 113824 153138 113876 153144
rect 114008 151904 114060 151910
rect 114008 151846 114060 151852
rect 114020 149954 114048 151846
rect 114296 149954 114324 171106
rect 114928 155508 114980 155514
rect 114928 155450 114980 155456
rect 114836 152516 114888 152522
rect 114836 152458 114888 152464
rect 114848 149954 114876 152458
rect 114940 150226 114968 155450
rect 115020 151836 115072 151842
rect 115124 151814 115152 527138
rect 116492 494080 116544 494086
rect 116492 494022 116544 494028
rect 115204 360256 115256 360262
rect 115204 360198 115256 360204
rect 115216 153134 115244 360198
rect 116504 161474 116532 494022
rect 116768 476196 116820 476202
rect 116768 476138 116820 476144
rect 116584 209840 116636 209846
rect 116584 209782 116636 209788
rect 116228 161446 116532 161474
rect 115204 153128 115256 153134
rect 115204 153070 115256 153076
rect 115848 152312 115900 152318
rect 115848 152254 115900 152260
rect 115124 151786 115428 151814
rect 115020 151778 115072 151784
rect 115032 150498 115060 151778
rect 115032 150470 115152 150498
rect 114940 150198 115014 150226
rect 113744 149926 113896 149954
rect 114020 149926 114172 149954
rect 114296 149926 114448 149954
rect 114724 149926 114876 149954
rect 114986 149940 115014 150198
rect 115124 149954 115152 150470
rect 115400 149954 115428 151786
rect 115860 149954 115888 152254
rect 116228 149954 116256 161446
rect 116492 158772 116544 158778
rect 116492 158714 116544 158720
rect 116308 153196 116360 153202
rect 116308 153138 116360 153144
rect 116320 150226 116348 153138
rect 116504 152998 116532 158714
rect 116596 153066 116624 209782
rect 116584 153060 116636 153066
rect 116584 153002 116636 153008
rect 116492 152992 116544 152998
rect 116492 152934 116544 152940
rect 116320 150198 116394 150226
rect 115124 149926 115276 149954
rect 115400 149926 115552 149954
rect 115828 149926 115888 149954
rect 116104 149926 116256 149954
rect 116366 149940 116394 150198
rect 116780 149954 116808 476138
rect 117044 443012 117096 443018
rect 117044 442954 117096 442960
rect 116952 151836 117004 151842
rect 116952 151778 117004 151784
rect 116964 149954 116992 151778
rect 116656 149926 116808 149954
rect 116932 149926 116992 149954
rect 117056 149954 117084 442954
rect 117596 426488 117648 426494
rect 117596 426430 117648 426436
rect 117504 155916 117556 155922
rect 117504 155858 117556 155864
rect 117516 149954 117544 155858
rect 117056 149926 117208 149954
rect 117484 149926 117544 149954
rect 117608 149954 117636 426430
rect 117872 393372 117924 393378
rect 117872 393314 117924 393320
rect 117780 152176 117832 152182
rect 117780 152118 117832 152124
rect 117792 151910 117820 152118
rect 117780 151904 117832 151910
rect 117780 151846 117832 151852
rect 117884 151814 117912 393314
rect 117964 376780 118016 376786
rect 117964 376722 118016 376728
rect 117976 154562 118004 376722
rect 118056 325712 118108 325718
rect 118056 325654 118108 325660
rect 118068 155922 118096 325654
rect 118148 226432 118200 226438
rect 118148 226374 118200 226380
rect 118056 155916 118108 155922
rect 118056 155858 118108 155864
rect 117964 154556 118016 154562
rect 117964 154498 118016 154504
rect 118160 153202 118188 226374
rect 118712 171134 118740 702406
rect 119344 342304 119396 342310
rect 119344 342246 119396 342252
rect 118712 171106 118832 171134
rect 118700 154556 118752 154562
rect 118700 154498 118752 154504
rect 118148 153196 118200 153202
rect 118148 153138 118200 153144
rect 118424 153128 118476 153134
rect 118424 153070 118476 153076
rect 118056 152516 118108 152522
rect 118056 152458 118108 152464
rect 118068 152250 118096 152458
rect 118056 152244 118108 152250
rect 118056 152186 118108 152192
rect 117884 151786 118188 151814
rect 118160 149954 118188 151786
rect 118436 149954 118464 153070
rect 118712 149954 118740 154498
rect 118804 154290 118832 171106
rect 118792 154284 118844 154290
rect 118792 154226 118844 154232
rect 119158 151872 119214 151881
rect 119158 151807 119214 151816
rect 119172 149954 119200 151807
rect 119356 150226 119384 342246
rect 119620 309188 119672 309194
rect 119620 309130 119672 309136
rect 119632 150226 119660 309130
rect 120632 292596 120684 292602
rect 120632 292538 120684 292544
rect 120448 259480 120500 259486
rect 120448 259422 120500 259428
rect 120356 242956 120408 242962
rect 120356 242898 120408 242904
rect 120368 156874 120396 242898
rect 120356 156868 120408 156874
rect 120356 156810 120408 156816
rect 120356 156596 120408 156602
rect 120356 156538 120408 156544
rect 119804 155916 119856 155922
rect 119804 155858 119856 155864
rect 119356 150198 119430 150226
rect 119632 150198 119706 150226
rect 117608 149926 117760 149954
rect 118160 149926 118312 149954
rect 118436 149926 118588 149954
rect 118712 149926 118864 149954
rect 119140 149926 119200 149954
rect 119402 149940 119430 150198
rect 119678 149940 119706 150198
rect 119816 149954 119844 155858
rect 120368 149954 120396 156538
rect 120460 150226 120488 259422
rect 120644 156602 120672 292538
rect 120724 276072 120776 276078
rect 120724 276014 120776 276020
rect 120632 156596 120684 156602
rect 120632 156538 120684 156544
rect 120736 150226 120764 276014
rect 121736 191888 121788 191894
rect 121736 191830 121788 191836
rect 120908 156868 120960 156874
rect 120908 156810 120960 156816
rect 120460 150198 120534 150226
rect 120736 150198 120810 150226
rect 119816 149926 119968 149954
rect 120244 149926 120396 149954
rect 120506 149940 120534 150198
rect 120782 149940 120810 150198
rect 120920 149954 120948 156810
rect 121460 153196 121512 153202
rect 121460 153138 121512 153144
rect 121184 153060 121236 153066
rect 121184 153002 121236 153008
rect 121196 149954 121224 153002
rect 121472 149954 121500 153138
rect 121748 149954 121776 191830
rect 122012 175296 122064 175302
rect 122012 175238 122064 175244
rect 122024 171134 122052 175238
rect 122024 171106 122328 171134
rect 122012 152992 122064 152998
rect 122012 152934 122064 152940
rect 122024 149954 122052 152934
rect 122300 149954 122328 171106
rect 139412 157078 139440 703582
rect 140424 703474 140452 703582
rect 140566 703520 140678 704960
rect 162186 703520 162298 704960
rect 183806 703520 183918 704960
rect 205426 703520 205538 704960
rect 227046 703520 227158 704960
rect 248666 703520 248778 704960
rect 269132 703582 270172 703610
rect 140608 703474 140636 703520
rect 140424 703446 140636 703474
rect 162228 700738 162256 703520
rect 183848 702434 183876 703520
rect 205468 703050 205496 703520
rect 204260 703044 204312 703050
rect 204260 702986 204312 702992
rect 205456 703044 205508 703050
rect 205456 702986 205508 702992
rect 183572 702406 183876 702434
rect 162216 700732 162268 700738
rect 162216 700674 162268 700680
rect 139400 157072 139452 157078
rect 139400 157014 139452 157020
rect 183572 155650 183600 702406
rect 204272 156942 204300 702986
rect 227088 700602 227116 703520
rect 248708 702434 248736 703520
rect 248432 702406 248736 702434
rect 227076 700596 227128 700602
rect 227076 700538 227128 700544
rect 204260 156936 204312 156942
rect 204260 156878 204312 156884
rect 183560 155644 183612 155650
rect 183560 155586 183612 155592
rect 248432 155446 248460 702406
rect 269132 156806 269160 703582
rect 270144 703474 270172 703582
rect 270286 703520 270398 704960
rect 291906 703520 292018 704960
rect 313526 703520 313638 704960
rect 335146 703520 335258 704960
rect 356072 703582 356652 703610
rect 270328 703474 270356 703520
rect 270144 703446 270356 703474
rect 291948 700534 291976 703520
rect 313568 702434 313596 703520
rect 335188 703050 335216 703520
rect 333980 703044 334032 703050
rect 333980 702986 334032 702992
rect 335176 703044 335228 703050
rect 335176 702986 335228 702992
rect 313292 702406 313596 702434
rect 291936 700528 291988 700534
rect 291936 700470 291988 700476
rect 269120 156800 269172 156806
rect 269120 156742 269172 156748
rect 248420 155440 248472 155446
rect 248420 155382 248472 155388
rect 313292 154154 313320 702406
rect 333992 156738 334020 702986
rect 333980 156732 334032 156738
rect 333980 156674 334032 156680
rect 356072 156670 356100 703582
rect 356624 703474 356652 703582
rect 356766 703520 356878 704960
rect 378386 703520 378498 704960
rect 398852 703582 399892 703610
rect 356808 703474 356836 703520
rect 356624 703446 356836 703474
rect 378428 702434 378456 703520
rect 378152 702406 378456 702434
rect 356060 156664 356112 156670
rect 356060 156606 356112 156612
rect 313280 154148 313332 154154
rect 313280 154090 313332 154096
rect 378152 154086 378180 702406
rect 398852 155378 398880 703582
rect 399864 703474 399892 703582
rect 400006 703520 400118 704960
rect 421626 703520 421738 704960
rect 443246 703520 443358 704960
rect 464866 703520 464978 704960
rect 486486 703520 486598 704960
rect 508106 703520 508218 704960
rect 528572 703582 529612 703610
rect 400048 703474 400076 703520
rect 399864 703446 400076 703474
rect 421668 700466 421696 703520
rect 443288 702434 443316 703520
rect 464908 703050 464936 703520
rect 463700 703044 463752 703050
rect 463700 702986 463752 702992
rect 464896 703044 464948 703050
rect 464896 702986 464948 702992
rect 443012 702406 443316 702434
rect 421656 700460 421708 700466
rect 421656 700402 421708 700408
rect 398840 155372 398892 155378
rect 398840 155314 398892 155320
rect 378140 154080 378192 154086
rect 378140 154022 378192 154028
rect 443012 154018 443040 702406
rect 463712 155310 463740 702986
rect 486528 700398 486556 703520
rect 508148 702434 508176 703520
rect 507872 702406 508176 702434
rect 486516 700392 486568 700398
rect 486516 700334 486568 700340
rect 463700 155304 463752 155310
rect 463700 155246 463752 155252
rect 443000 154012 443052 154018
rect 443000 153954 443052 153960
rect 507872 153950 507900 702406
rect 528572 155242 528600 703582
rect 529584 703474 529612 703582
rect 529726 703520 529838 704960
rect 551346 703520 551458 704960
rect 572966 703520 573078 704960
rect 529768 703474 529796 703520
rect 529584 703446 529796 703474
rect 551388 700330 551416 703520
rect 573008 702434 573036 703520
rect 572732 702406 573036 702434
rect 551376 700324 551428 700330
rect 551376 700266 551428 700272
rect 528560 155236 528612 155242
rect 528560 155178 528612 155184
rect 507860 153944 507912 153950
rect 507860 153886 507912 153892
rect 572732 153882 572760 702406
rect 580170 696008 580226 696017
rect 580170 695943 580226 695952
rect 580184 695570 580212 695943
rect 580172 695564 580224 695570
rect 580172 695506 580224 695512
rect 580172 680400 580224 680406
rect 580170 680368 580172 680377
rect 580224 680368 580226 680377
rect 580170 680303 580226 680312
rect 580170 664728 580226 664737
rect 580170 664663 580226 664672
rect 580184 663814 580212 664663
rect 580172 663808 580224 663814
rect 580172 663750 580224 663756
rect 580170 649088 580226 649097
rect 580170 649023 580226 649032
rect 580184 648650 580212 649023
rect 580172 648644 580224 648650
rect 580172 648586 580224 648592
rect 580172 633480 580224 633486
rect 580170 633448 580172 633457
rect 580224 633448 580226 633457
rect 580170 633383 580226 633392
rect 580170 617808 580226 617817
rect 580170 617743 580226 617752
rect 580184 616894 580212 617743
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 602168 580226 602177
rect 580170 602103 580226 602112
rect 580184 601730 580212 602103
rect 580172 601724 580224 601730
rect 580172 601666 580224 601672
rect 580908 586560 580960 586566
rect 580906 586528 580908 586537
rect 580960 586528 580962 586537
rect 580906 586463 580962 586472
rect 580170 570888 580226 570897
rect 580170 570823 580226 570832
rect 580184 569974 580212 570823
rect 580172 569968 580224 569974
rect 580172 569910 580224 569916
rect 580170 555248 580226 555257
rect 580170 555183 580226 555192
rect 580184 554810 580212 555183
rect 580172 554804 580224 554810
rect 580172 554746 580224 554752
rect 580172 539640 580224 539646
rect 580170 539608 580172 539617
rect 580224 539608 580226 539617
rect 580170 539543 580226 539552
rect 580170 523968 580226 523977
rect 580170 523903 580226 523912
rect 580184 523054 580212 523903
rect 580172 523048 580224 523054
rect 580172 522990 580224 522996
rect 580170 508328 580226 508337
rect 580170 508263 580226 508272
rect 580184 507890 580212 508263
rect 580172 507884 580224 507890
rect 580172 507826 580224 507832
rect 580172 492720 580224 492726
rect 580170 492688 580172 492697
rect 580224 492688 580226 492697
rect 580170 492623 580226 492632
rect 580170 477048 580226 477057
rect 580170 476983 580226 476992
rect 580184 476134 580212 476983
rect 580172 476128 580224 476134
rect 580172 476070 580224 476076
rect 580170 461408 580226 461417
rect 580170 461343 580226 461352
rect 580184 460970 580212 461343
rect 580172 460964 580224 460970
rect 580172 460906 580224 460912
rect 580172 445800 580224 445806
rect 580170 445768 580172 445777
rect 580224 445768 580226 445777
rect 580170 445703 580226 445712
rect 580170 430128 580226 430137
rect 580170 430063 580226 430072
rect 580184 429214 580212 430063
rect 580172 429208 580224 429214
rect 580172 429150 580224 429156
rect 580170 414488 580226 414497
rect 580170 414423 580226 414432
rect 580184 414050 580212 414423
rect 580172 414044 580224 414050
rect 580172 413986 580224 413992
rect 580172 398880 580224 398886
rect 580170 398848 580172 398857
rect 580224 398848 580226 398857
rect 580170 398783 580226 398792
rect 580170 383208 580226 383217
rect 580170 383143 580226 383152
rect 580184 382294 580212 383143
rect 580172 382288 580224 382294
rect 580172 382230 580224 382236
rect 580170 367568 580226 367577
rect 580170 367503 580226 367512
rect 580184 367130 580212 367503
rect 580172 367124 580224 367130
rect 580172 367066 580224 367072
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 336288 580226 336297
rect 580170 336223 580226 336232
rect 580184 335374 580212 336223
rect 580172 335368 580224 335374
rect 580172 335310 580224 335316
rect 580170 320648 580226 320657
rect 580170 320583 580226 320592
rect 580184 320210 580212 320583
rect 580172 320204 580224 320210
rect 580172 320146 580224 320152
rect 580172 305040 580224 305046
rect 580170 305008 580172 305017
rect 580224 305008 580226 305017
rect 580170 304943 580226 304952
rect 580170 289368 580226 289377
rect 580170 289303 580226 289312
rect 580184 288454 580212 289303
rect 580172 288448 580224 288454
rect 580172 288390 580224 288396
rect 580170 273728 580226 273737
rect 580170 273663 580226 273672
rect 580184 273290 580212 273663
rect 580172 273284 580224 273290
rect 580172 273226 580224 273232
rect 580908 258120 580960 258126
rect 580906 258088 580908 258097
rect 580960 258088 580962 258097
rect 580906 258023 580962 258032
rect 580170 242448 580226 242457
rect 580170 242383 580226 242392
rect 580184 241534 580212 242383
rect 580172 241528 580224 241534
rect 580172 241470 580224 241476
rect 580170 226808 580226 226817
rect 580170 226743 580226 226752
rect 580184 226370 580212 226743
rect 580172 226364 580224 226370
rect 580172 226306 580224 226312
rect 580172 211200 580224 211206
rect 580170 211168 580172 211177
rect 580224 211168 580226 211177
rect 580170 211103 580226 211112
rect 580170 195528 580226 195537
rect 580170 195463 580226 195472
rect 580184 194614 580212 195463
rect 580172 194608 580224 194614
rect 580172 194550 580224 194556
rect 580170 179888 580226 179897
rect 580170 179823 580226 179832
rect 580184 179450 580212 179823
rect 580172 179444 580224 179450
rect 580172 179386 580224 179392
rect 580172 164280 580224 164286
rect 580170 164248 580172 164257
rect 580224 164248 580226 164257
rect 580170 164183 580226 164192
rect 572720 153876 572772 153882
rect 572720 153818 572772 153824
rect 128728 152924 128780 152930
rect 128728 152866 128780 152872
rect 123116 152856 123168 152862
rect 123116 152798 123168 152804
rect 122840 152720 122892 152726
rect 122840 152662 122892 152668
rect 122852 149954 122880 152662
rect 123128 149954 123156 152798
rect 123944 152380 123996 152386
rect 123944 152322 123996 152328
rect 123392 150748 123444 150754
rect 123392 150690 123444 150696
rect 123404 149954 123432 150690
rect 123668 150680 123720 150686
rect 123668 150622 123720 150628
rect 123680 149954 123708 150622
rect 123956 149954 123984 152322
rect 127992 152312 128044 152318
rect 127992 152254 128044 152260
rect 124770 152144 124826 152153
rect 124770 152079 124826 152088
rect 124220 150612 124272 150618
rect 124220 150554 124272 150560
rect 124232 149954 124260 150554
rect 124496 150544 124548 150550
rect 124496 150486 124548 150492
rect 124508 149954 124536 150486
rect 124784 149954 124812 152079
rect 120920 149926 121072 149954
rect 121196 149926 121348 149954
rect 121472 149926 121624 149954
rect 121748 149926 121900 149954
rect 122024 149926 122176 149954
rect 122300 149926 122452 149954
rect 122852 149926 123004 149954
rect 123128 149926 123280 149954
rect 123404 149926 123556 149954
rect 123680 149926 123832 149954
rect 123956 149926 124108 149954
rect 124232 149926 124384 149954
rect 124508 149926 124660 149954
rect 124784 149926 124936 149954
rect 93584 149864 93636 149870
rect 90284 149802 90436 149818
rect 112352 149864 112404 149870
rect 93636 149812 93748 149818
rect 93584 149806 93748 149812
rect 112352 149806 112404 149812
rect 112628 149864 112680 149870
rect 112680 149812 112792 149818
rect 112628 149806 112792 149812
rect 90272 149796 90436 149802
rect 90324 149790 90436 149796
rect 93596 149790 93748 149806
rect 112640 149790 112792 149806
rect 90272 149738 90324 149744
rect 89168 149728 89220 149734
rect 85192 149666 85344 149682
rect 92480 149728 92532 149734
rect 89220 149676 89332 149682
rect 89168 149670 89332 149676
rect 92532 149676 92644 149682
rect 92480 149670 92644 149676
rect 85192 149660 85356 149666
rect 85192 149654 85304 149660
rect 89180 149654 89332 149670
rect 89444 149660 89496 149666
rect 85304 149602 85356 149608
rect 89444 149602 89496 149608
rect 91652 149660 91704 149666
rect 92492 149654 92644 149670
rect 91652 149602 91704 149608
rect 86960 149592 87012 149598
rect 85868 149530 86020 149546
rect 85856 149524 86020 149530
rect 85908 149518 86020 149524
rect 86572 149530 86724 149546
rect 87510 149560 87566 149569
rect 87012 149540 87124 149546
rect 86960 149534 87124 149540
rect 86572 149524 86736 149530
rect 86572 149518 86684 149524
rect 85856 149466 85908 149472
rect 86972 149518 87124 149534
rect 87400 149518 87510 149546
rect 87510 149495 87566 149504
rect 86684 149466 86736 149472
rect 89456 149462 89484 149602
rect 91664 149462 91692 149602
rect 91928 149592 91980 149598
rect 118148 149592 118200 149598
rect 91928 149534 91980 149540
rect 94134 149560 94190 149569
rect 91940 149462 91968 149534
rect 118036 149540 118148 149546
rect 118036 149534 118200 149540
rect 118036 149518 118188 149534
rect 94134 149495 94190 149504
rect 94148 149462 94176 149495
rect 84568 149456 84620 149462
rect 86408 149456 86460 149462
rect 84620 149404 84916 149410
rect 84568 149398 84916 149404
rect 84580 149382 84916 149398
rect 86296 149404 86408 149410
rect 89444 149456 89496 149462
rect 86296 149398 86460 149404
rect 88062 149424 88118 149433
rect 86296 149382 86448 149398
rect 88118 149382 88228 149410
rect 89444 149398 89496 149404
rect 91652 149456 91704 149462
rect 91652 149398 91704 149404
rect 91928 149456 91980 149462
rect 91928 149398 91980 149404
rect 94136 149456 94188 149462
rect 94136 149398 94188 149404
rect 122564 149456 122616 149462
rect 122616 149404 122728 149410
rect 122564 149398 122728 149404
rect 122576 149382 122728 149398
rect 88062 149359 88118 149368
rect 82360 101516 82412 101522
rect 82360 101458 82412 101464
rect 97586 100224 97638 100230
rect 97586 100166 97638 100172
rect 97598 100164 97626 100166
rect 86650 100162 86678 100164
rect 98978 100162 99006 100164
rect 117654 100162 117682 100164
rect 121610 100162 121638 100164
rect 128004 100162 128032 152254
rect 128544 152244 128596 152250
rect 128544 152186 128596 152192
rect 128452 152176 128504 152182
rect 128452 152118 128504 152124
rect 128360 152108 128412 152114
rect 128360 152050 128412 152056
rect 128176 151836 128228 151842
rect 128176 151778 128228 151784
rect 128084 149592 128136 149598
rect 128084 149534 128136 149540
rect 86638 100156 86690 100162
rect 86638 100098 86690 100104
rect 98966 100156 99018 100162
rect 98966 100098 99018 100104
rect 117642 100156 117694 100162
rect 117642 100098 117694 100104
rect 121598 100156 121650 100162
rect 121598 100098 121650 100104
rect 127992 100156 128044 100162
rect 127992 100098 128044 100104
rect 90502 100088 90554 100094
rect 90502 100030 90554 100036
rect 93722 100088 93774 100094
rect 93722 100030 93774 100036
rect 99610 100088 99662 100094
rect 99610 100030 99662 100036
rect 100714 100088 100766 100094
rect 100714 100030 100766 100036
rect 104854 100088 104906 100094
rect 104854 100030 104906 100036
rect 107338 100088 107390 100094
rect 107338 100030 107390 100036
rect 112582 100088 112634 100094
rect 112582 100030 112634 100036
rect 121322 100088 121374 100094
rect 121322 100030 121374 100036
rect 125738 100088 125790 100094
rect 125738 100030 125790 100036
rect 127118 100088 127170 100094
rect 127808 100088 127860 100094
rect 127118 100030 127170 100036
rect 90514 100028 90542 100030
rect 93734 100028 93762 100030
rect 99622 100028 99650 100030
rect 100726 100028 100754 100030
rect 104866 100028 104894 100030
rect 107350 100028 107378 100030
rect 112594 100028 112622 100030
rect 121334 100028 121362 100030
rect 125750 100028 125778 100030
rect 127130 100028 127158 100030
rect 82360 99952 82412 99958
rect 82360 99894 82412 99900
rect 82268 96552 82320 96558
rect 82268 96494 82320 96500
rect 82372 96218 82400 99894
rect 82510 99770 82538 100028
rect 82602 99890 82630 100028
rect 82590 99884 82642 99890
rect 82590 99826 82642 99832
rect 82694 99770 82722 100028
rect 82786 99890 82814 100028
rect 82774 99884 82826 99890
rect 82774 99826 82826 99832
rect 82878 99770 82906 100028
rect 82464 99742 82538 99770
rect 82648 99742 82722 99770
rect 82832 99742 82906 99770
rect 82970 99770 82998 100028
rect 83062 99890 83090 100028
rect 83050 99884 83102 99890
rect 83050 99826 83102 99832
rect 83154 99770 83182 100028
rect 83246 99822 83274 100028
rect 83338 99890 83366 100028
rect 83326 99884 83378 99890
rect 83326 99826 83378 99832
rect 82970 99742 83044 99770
rect 82360 96212 82412 96218
rect 82360 96154 82412 96160
rect 82464 94722 82492 99742
rect 82648 99374 82676 99742
rect 82556 99346 82676 99374
rect 82452 94716 82504 94722
rect 82452 94658 82504 94664
rect 82556 94568 82584 99346
rect 82728 98320 82780 98326
rect 82728 98262 82780 98268
rect 82636 96688 82688 96694
rect 82636 96630 82688 96636
rect 82464 94540 82584 94568
rect 82464 4962 82492 94540
rect 82648 94500 82676 96630
rect 82556 94472 82676 94500
rect 82556 44878 82584 94472
rect 82740 89714 82768 98262
rect 82832 97306 82860 99742
rect 82912 99680 82964 99686
rect 82912 99622 82964 99628
rect 82820 97300 82872 97306
rect 82820 97242 82872 97248
rect 82924 94450 82952 99622
rect 82912 94444 82964 94450
rect 82912 94386 82964 94392
rect 82648 89686 82768 89714
rect 82648 45014 82676 89686
rect 82636 45008 82688 45014
rect 82636 44950 82688 44956
rect 82544 44872 82596 44878
rect 82544 44814 82596 44820
rect 82452 4956 82504 4962
rect 82452 4898 82504 4904
rect 82360 4820 82412 4826
rect 82360 4762 82412 4768
rect 82372 2854 82400 4762
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 82360 2848 82412 2854
rect 82360 2790 82412 2796
rect 82740 480 82768 3470
rect 83016 3466 83044 99742
rect 83108 99742 83182 99770
rect 83234 99816 83286 99822
rect 83430 99770 83458 100028
rect 83522 99958 83550 100028
rect 83614 99958 83642 100028
rect 83510 99952 83562 99958
rect 83510 99894 83562 99900
rect 83602 99952 83654 99958
rect 83706 99929 83734 100028
rect 83602 99894 83654 99900
rect 83692 99920 83748 99929
rect 83692 99855 83748 99864
rect 83798 99822 83826 100028
rect 83234 99758 83286 99764
rect 83384 99742 83458 99770
rect 83786 99816 83838 99822
rect 83786 99758 83838 99764
rect 83108 96694 83136 99742
rect 83188 99680 83240 99686
rect 83384 99634 83412 99742
rect 83188 99622 83240 99628
rect 83096 96688 83148 96694
rect 83096 96630 83148 96636
rect 83096 94580 83148 94586
rect 83096 94522 83148 94528
rect 83108 3670 83136 94522
rect 83200 5302 83228 99622
rect 83292 99606 83412 99634
rect 83556 99680 83608 99686
rect 83556 99622 83608 99628
rect 83648 99680 83700 99686
rect 83890 99668 83918 100028
rect 83982 99770 84010 100028
rect 84074 99958 84102 100028
rect 84166 99958 84194 100028
rect 84258 99958 84286 100028
rect 84350 99958 84378 100028
rect 84062 99952 84114 99958
rect 84062 99894 84114 99900
rect 84154 99952 84206 99958
rect 84154 99894 84206 99900
rect 84246 99952 84298 99958
rect 84246 99894 84298 99900
rect 84338 99952 84390 99958
rect 84442 99929 84470 100028
rect 84338 99894 84390 99900
rect 84428 99920 84484 99929
rect 84428 99855 84484 99864
rect 84384 99816 84436 99822
rect 84290 99784 84346 99793
rect 83982 99742 84056 99770
rect 83648 99622 83700 99628
rect 83752 99640 83918 99668
rect 83292 6186 83320 99606
rect 83372 99544 83424 99550
rect 83372 99486 83424 99492
rect 83384 98190 83412 99486
rect 83462 99388 83518 99397
rect 83462 99323 83518 99332
rect 83372 98184 83424 98190
rect 83372 98126 83424 98132
rect 83372 94716 83424 94722
rect 83372 94658 83424 94664
rect 83384 6254 83412 94658
rect 83476 94586 83504 99323
rect 83464 94580 83516 94586
rect 83464 94522 83516 94528
rect 83568 94450 83596 99622
rect 83660 94722 83688 99622
rect 83648 94716 83700 94722
rect 83648 94658 83700 94664
rect 83752 94568 83780 99640
rect 83832 99544 83884 99550
rect 83832 99486 83884 99492
rect 83660 94540 83780 94568
rect 83464 94444 83516 94450
rect 83464 94386 83516 94392
rect 83556 94444 83608 94450
rect 83556 94386 83608 94392
rect 83476 7614 83504 94386
rect 83556 84244 83608 84250
rect 83556 84186 83608 84192
rect 83568 16574 83596 84186
rect 83660 21418 83688 94540
rect 83740 94444 83792 94450
rect 83740 94386 83792 94392
rect 83648 21412 83700 21418
rect 83648 21354 83700 21360
rect 83568 16546 83688 16574
rect 83464 7608 83516 7614
rect 83464 7550 83516 7556
rect 83372 6248 83424 6254
rect 83372 6190 83424 6196
rect 83280 6180 83332 6186
rect 83280 6122 83332 6128
rect 83188 5296 83240 5302
rect 83188 5238 83240 5244
rect 83096 3664 83148 3670
rect 83096 3606 83148 3612
rect 83660 3482 83688 16546
rect 83752 4146 83780 94386
rect 83844 16574 83872 99486
rect 83924 98184 83976 98190
rect 83924 98126 83976 98132
rect 83936 84930 83964 98126
rect 84028 87650 84056 99742
rect 84200 99748 84252 99754
rect 84534 99770 84562 100028
rect 84626 99890 84654 100028
rect 84718 99890 84746 100028
rect 84614 99884 84666 99890
rect 84614 99826 84666 99832
rect 84706 99884 84758 99890
rect 84706 99826 84758 99832
rect 84810 99770 84838 100028
rect 84902 99793 84930 100028
rect 84384 99758 84436 99764
rect 84290 99719 84346 99728
rect 84200 99690 84252 99696
rect 84212 98297 84240 99690
rect 84198 98288 84254 98297
rect 84198 98223 84254 98232
rect 84304 97646 84332 99719
rect 84292 97640 84344 97646
rect 84292 97582 84344 97588
rect 84396 97578 84424 99758
rect 84488 99742 84562 99770
rect 84764 99742 84838 99770
rect 84888 99784 84944 99793
rect 84488 99686 84516 99742
rect 84476 99680 84528 99686
rect 84476 99622 84528 99628
rect 84476 99544 84528 99550
rect 84476 99486 84528 99492
rect 84384 97572 84436 97578
rect 84384 97514 84436 97520
rect 84384 97436 84436 97442
rect 84384 97378 84436 97384
rect 84396 94382 84424 97378
rect 84384 94376 84436 94382
rect 84384 94318 84436 94324
rect 84016 87644 84068 87650
rect 84016 87586 84068 87592
rect 83924 84924 83976 84930
rect 83924 84866 83976 84872
rect 83844 16546 83964 16574
rect 83740 4140 83792 4146
rect 83740 4082 83792 4088
rect 83936 3738 83964 16546
rect 84488 5030 84516 99486
rect 84568 99476 84620 99482
rect 84568 99418 84620 99424
rect 84660 99476 84712 99482
rect 84660 99418 84712 99424
rect 84580 6322 84608 99418
rect 84672 6390 84700 99418
rect 84764 94790 84792 99742
rect 84888 99719 84944 99728
rect 84994 99668 85022 100028
rect 85086 99929 85114 100028
rect 85178 99958 85206 100028
rect 85166 99952 85218 99958
rect 85072 99920 85128 99929
rect 85166 99894 85218 99900
rect 85072 99855 85128 99864
rect 85270 99770 85298 100028
rect 85362 99822 85390 100028
rect 85224 99742 85298 99770
rect 85350 99816 85402 99822
rect 85350 99758 85402 99764
rect 85454 99770 85482 100028
rect 85546 99929 85574 100028
rect 85532 99920 85588 99929
rect 85532 99855 85588 99864
rect 85638 99822 85666 100028
rect 85730 99929 85758 100028
rect 85716 99920 85772 99929
rect 85822 99890 85850 100028
rect 85914 99890 85942 100028
rect 86006 99958 86034 100028
rect 85994 99952 86046 99958
rect 85994 99894 86046 99900
rect 85716 99855 85772 99864
rect 85810 99884 85862 99890
rect 85810 99826 85862 99832
rect 85902 99884 85954 99890
rect 85902 99826 85954 99832
rect 85626 99816 85678 99822
rect 85454 99742 85528 99770
rect 86098 99804 86126 100028
rect 86190 99958 86218 100028
rect 86282 99958 86310 100028
rect 86178 99952 86230 99958
rect 86178 99894 86230 99900
rect 86270 99952 86322 99958
rect 86374 99929 86402 100028
rect 86270 99894 86322 99900
rect 86360 99920 86416 99929
rect 86360 99855 86416 99864
rect 86466 99822 86494 100028
rect 86558 99906 86586 100028
rect 86558 99890 86632 99906
rect 86558 99884 86644 99890
rect 86558 99878 86592 99884
rect 86592 99826 86644 99832
rect 86742 99822 86770 100028
rect 86834 99929 86862 100028
rect 86820 99920 86876 99929
rect 86820 99855 86876 99864
rect 86316 99816 86368 99822
rect 85626 99758 85678 99764
rect 85762 99784 85818 99793
rect 84994 99640 85068 99668
rect 84936 99476 84988 99482
rect 84936 99418 84988 99424
rect 84844 99408 84896 99414
rect 84844 99350 84896 99356
rect 84752 94784 84804 94790
rect 84752 94726 84804 94732
rect 84856 94568 84884 99350
rect 84764 94540 84884 94568
rect 84948 94568 84976 99418
rect 85040 94722 85068 99640
rect 85224 99482 85252 99742
rect 85396 99680 85448 99686
rect 85396 99622 85448 99628
rect 85304 99612 85356 99618
rect 85304 99554 85356 99560
rect 85212 99476 85264 99482
rect 85212 99418 85264 99424
rect 85210 99376 85266 99385
rect 85210 99311 85266 99320
rect 85120 94784 85172 94790
rect 85120 94726 85172 94732
rect 85028 94716 85080 94722
rect 85028 94658 85080 94664
rect 84948 94540 85068 94568
rect 84764 44946 84792 94540
rect 84844 94444 84896 94450
rect 84844 94386 84896 94392
rect 84752 44940 84804 44946
rect 84752 44882 84804 44888
rect 84752 20052 84804 20058
rect 84752 19994 84804 20000
rect 84660 6384 84712 6390
rect 84660 6326 84712 6332
rect 84568 6316 84620 6322
rect 84568 6258 84620 6264
rect 84476 5024 84528 5030
rect 84476 4966 84528 4972
rect 83924 3732 83976 3738
rect 83924 3674 83976 3680
rect 84764 3482 84792 19994
rect 84856 6458 84884 94386
rect 84936 94376 84988 94382
rect 84936 94318 84988 94324
rect 84948 6730 84976 94318
rect 84936 6724 84988 6730
rect 84936 6666 84988 6672
rect 84844 6452 84896 6458
rect 84844 6394 84896 6400
rect 85040 5234 85068 94540
rect 85028 5228 85080 5234
rect 85028 5170 85080 5176
rect 85132 5098 85160 94726
rect 85224 86290 85252 99311
rect 85316 94450 85344 99554
rect 85408 96614 85436 99622
rect 85500 97034 85528 99742
rect 86098 99776 86172 99804
rect 85762 99719 85818 99728
rect 85672 99680 85724 99686
rect 85672 99622 85724 99628
rect 85776 99634 85804 99719
rect 86040 99680 86092 99686
rect 85946 99648 86002 99657
rect 85684 98297 85712 99622
rect 85776 99606 85896 99634
rect 85670 98288 85726 98297
rect 85670 98223 85726 98232
rect 85764 97504 85816 97510
rect 85764 97446 85816 97452
rect 85488 97028 85540 97034
rect 85488 96970 85540 96976
rect 85672 96620 85724 96626
rect 85408 96586 85528 96614
rect 85396 94716 85448 94722
rect 85396 94658 85448 94664
rect 85304 94444 85356 94450
rect 85304 94386 85356 94392
rect 85212 86284 85264 86290
rect 85212 86226 85264 86232
rect 85408 5166 85436 94658
rect 85500 87718 85528 96586
rect 85672 96562 85724 96568
rect 85488 87712 85540 87718
rect 85488 87654 85540 87660
rect 85684 84194 85712 96562
rect 85592 84166 85712 84194
rect 85592 83502 85620 84166
rect 85580 83496 85632 83502
rect 85580 83438 85632 83444
rect 85396 5160 85448 5166
rect 85396 5102 85448 5108
rect 85120 5092 85172 5098
rect 85120 5034 85172 5040
rect 85776 3806 85804 97446
rect 85868 94586 85896 99606
rect 86040 99622 86092 99628
rect 85946 99583 86002 99592
rect 85856 94580 85908 94586
rect 85856 94522 85908 94528
rect 85960 94500 85988 99583
rect 86052 94568 86080 99622
rect 86144 97510 86172 99776
rect 86314 99784 86316 99793
rect 86454 99816 86506 99822
rect 86368 99784 86370 99793
rect 86454 99758 86506 99764
rect 86730 99816 86782 99822
rect 86730 99758 86782 99764
rect 86314 99719 86370 99728
rect 86592 99748 86644 99754
rect 86926 99736 86954 100028
rect 87018 99958 87046 100028
rect 87006 99952 87058 99958
rect 87006 99894 87058 99900
rect 87110 99804 87138 100028
rect 87202 99822 87230 100028
rect 87294 99822 87322 100028
rect 87064 99776 87138 99804
rect 87190 99816 87242 99822
rect 86926 99708 87000 99736
rect 86592 99690 86644 99696
rect 86408 99612 86460 99618
rect 86408 99554 86460 99560
rect 86224 99408 86276 99414
rect 86224 99350 86276 99356
rect 86132 97504 86184 97510
rect 86132 97446 86184 97452
rect 86052 94540 86172 94568
rect 85960 94472 86080 94500
rect 85856 94444 85908 94450
rect 85856 94386 85908 94392
rect 85868 5370 85896 94386
rect 85948 94376 86000 94382
rect 85948 94318 86000 94324
rect 85960 6798 85988 94318
rect 85948 6792 86000 6798
rect 85948 6734 86000 6740
rect 86052 6662 86080 94472
rect 86040 6656 86092 6662
rect 86040 6598 86092 6604
rect 86144 6526 86172 94540
rect 86236 6594 86264 99350
rect 86420 97442 86448 99554
rect 86604 98326 86632 99690
rect 86776 99680 86828 99686
rect 86776 99622 86828 99628
rect 86866 99648 86922 99657
rect 86684 99476 86736 99482
rect 86684 99418 86736 99424
rect 86592 98320 86644 98326
rect 86498 98288 86554 98297
rect 86592 98262 86644 98268
rect 86498 98223 86554 98232
rect 86408 97436 86460 97442
rect 86408 97378 86460 97384
rect 86408 96688 86460 96694
rect 86408 96630 86460 96636
rect 86316 94580 86368 94586
rect 86316 94522 86368 94528
rect 86328 7682 86356 94522
rect 86420 84250 86448 96630
rect 86512 89714 86540 98223
rect 86512 89686 86632 89714
rect 86408 84244 86460 84250
rect 86408 84186 86460 84192
rect 86316 7676 86368 7682
rect 86316 7618 86368 7624
rect 86224 6588 86276 6594
rect 86224 6530 86276 6536
rect 86132 6520 86184 6526
rect 86132 6462 86184 6468
rect 85856 5364 85908 5370
rect 85856 5306 85908 5312
rect 86604 3874 86632 89686
rect 86696 3942 86724 99418
rect 86788 94382 86816 99622
rect 86866 99583 86922 99592
rect 86880 94450 86908 99583
rect 86972 94586 87000 99708
rect 87064 99464 87092 99776
rect 87190 99758 87242 99764
rect 87282 99816 87334 99822
rect 87282 99758 87334 99764
rect 87386 99770 87414 100028
rect 87478 99929 87506 100028
rect 87464 99920 87520 99929
rect 87570 99890 87598 100028
rect 87464 99855 87520 99864
rect 87558 99884 87610 99890
rect 87558 99826 87610 99832
rect 87386 99742 87460 99770
rect 87432 99657 87460 99742
rect 87512 99748 87564 99754
rect 87512 99690 87564 99696
rect 87418 99648 87474 99657
rect 87144 99612 87196 99618
rect 87196 99572 87276 99600
rect 87418 99583 87474 99592
rect 87144 99554 87196 99560
rect 87064 99436 87184 99464
rect 87052 99340 87104 99346
rect 87052 99282 87104 99288
rect 86960 94580 87012 94586
rect 87064 94568 87092 99282
rect 87156 94722 87184 99436
rect 87248 94722 87276 99572
rect 87420 99544 87472 99550
rect 87326 99512 87382 99521
rect 87420 99486 87472 99492
rect 87326 99447 87382 99456
rect 87144 94716 87196 94722
rect 87144 94658 87196 94664
rect 87236 94716 87288 94722
rect 87236 94658 87288 94664
rect 87064 94540 87276 94568
rect 86960 94522 87012 94528
rect 86868 94444 86920 94450
rect 86868 94386 86920 94392
rect 87144 94444 87196 94450
rect 87144 94386 87196 94392
rect 86776 94376 86828 94382
rect 86776 94318 86828 94324
rect 86684 3936 86736 3942
rect 86684 3878 86736 3884
rect 86592 3868 86644 3874
rect 86592 3810 86644 3816
rect 85764 3800 85816 3806
rect 85764 3742 85816 3748
rect 86040 3528 86092 3534
rect 83004 3460 83056 3466
rect 83660 3454 83872 3482
rect 84764 3454 84976 3482
rect 86040 3470 86092 3476
rect 83004 3402 83056 3408
rect 83844 480 83872 3454
rect 84948 480 84976 3454
rect 86052 480 86080 3470
rect 87156 3194 87184 94386
rect 87248 3534 87276 94540
rect 87340 3602 87368 99447
rect 87432 96762 87460 99486
rect 87420 96756 87472 96762
rect 87420 96698 87472 96704
rect 87524 96694 87552 99690
rect 87662 99668 87690 100028
rect 87754 99770 87782 100028
rect 87846 99958 87874 100028
rect 87834 99952 87886 99958
rect 87834 99894 87886 99900
rect 87938 99804 87966 100028
rect 88030 99958 88058 100028
rect 88018 99952 88070 99958
rect 88122 99929 88150 100028
rect 88018 99894 88070 99900
rect 88108 99920 88164 99929
rect 88108 99855 88164 99864
rect 87938 99793 88104 99804
rect 87938 99784 88118 99793
rect 87938 99776 88062 99784
rect 87754 99742 87828 99770
rect 87662 99640 87736 99668
rect 87604 99544 87656 99550
rect 87604 99486 87656 99492
rect 87512 96688 87564 96694
rect 87512 96630 87564 96636
rect 87616 94738 87644 99486
rect 87708 95234 87736 99640
rect 87800 99618 87828 99742
rect 88214 99736 88242 100028
rect 88306 99890 88334 100028
rect 88294 99884 88346 99890
rect 88294 99826 88346 99832
rect 88398 99827 88426 100028
rect 88490 99958 88518 100028
rect 88582 99958 88610 100028
rect 88478 99952 88530 99958
rect 88478 99894 88530 99900
rect 88570 99952 88622 99958
rect 88570 99894 88622 99900
rect 88384 99818 88440 99827
rect 88384 99753 88440 99762
rect 88674 99736 88702 100028
rect 88766 99890 88794 100028
rect 88754 99884 88806 99890
rect 88754 99826 88806 99832
rect 88858 99770 88886 100028
rect 88950 99958 88978 100028
rect 88938 99952 88990 99958
rect 88938 99894 88990 99900
rect 89042 99770 89070 100028
rect 89134 99963 89162 100028
rect 89120 99954 89176 99963
rect 89226 99958 89254 100028
rect 89318 99958 89346 100028
rect 89120 99889 89176 99898
rect 89214 99952 89266 99958
rect 89214 99894 89266 99900
rect 89306 99952 89358 99958
rect 89306 99894 89358 99900
rect 89410 99804 89438 100028
rect 89502 99822 89530 100028
rect 89594 99958 89622 100028
rect 89582 99952 89634 99958
rect 89582 99894 89634 99900
rect 89364 99776 89438 99804
rect 89490 99816 89542 99822
rect 88858 99742 88932 99770
rect 89042 99742 89116 99770
rect 88062 99719 88118 99728
rect 88168 99708 88242 99736
rect 88628 99708 88702 99736
rect 87880 99680 87932 99686
rect 87932 99640 88012 99668
rect 87880 99622 87932 99628
rect 87788 99612 87840 99618
rect 87788 99554 87840 99560
rect 87880 99544 87932 99550
rect 87786 99512 87842 99521
rect 87880 99486 87932 99492
rect 87786 99447 87842 99456
rect 87800 97102 87828 99447
rect 87788 97096 87840 97102
rect 87788 97038 87840 97044
rect 87708 95206 87828 95234
rect 87512 94716 87564 94722
rect 87616 94710 87736 94738
rect 87512 94658 87564 94664
rect 87420 94512 87472 94518
rect 87420 94454 87472 94460
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 87236 3528 87288 3534
rect 87236 3470 87288 3476
rect 87432 3466 87460 94454
rect 87524 4078 87552 94658
rect 87604 94580 87656 94586
rect 87604 94522 87656 94528
rect 87512 4072 87564 4078
rect 87512 4014 87564 4020
rect 87616 4010 87644 94522
rect 87708 4826 87736 94710
rect 87800 20058 87828 95206
rect 87892 94450 87920 99486
rect 87880 94444 87932 94450
rect 87880 94386 87932 94392
rect 87788 20052 87840 20058
rect 87788 19994 87840 20000
rect 87984 6914 88012 99640
rect 88062 99648 88118 99657
rect 88168 99618 88196 99708
rect 88340 99680 88392 99686
rect 88340 99622 88392 99628
rect 88062 99583 88118 99592
rect 88156 99612 88208 99618
rect 88076 94518 88104 99583
rect 88156 99554 88208 99560
rect 88154 99512 88210 99521
rect 88154 99447 88210 99456
rect 88064 94512 88116 94518
rect 88064 94454 88116 94460
rect 88064 94376 88116 94382
rect 88064 94318 88116 94324
rect 88076 87786 88104 94318
rect 88064 87780 88116 87786
rect 88064 87722 88116 87728
rect 88168 16574 88196 99447
rect 88352 94586 88380 99622
rect 88522 99512 88578 99521
rect 88432 99476 88484 99482
rect 88522 99447 88578 99456
rect 88432 99418 88484 99424
rect 88444 97730 88472 99418
rect 88536 98376 88564 99447
rect 88628 98530 88656 99708
rect 88904 99634 88932 99742
rect 88812 99606 88932 99634
rect 88984 99680 89036 99686
rect 88984 99622 89036 99628
rect 89088 99634 89116 99742
rect 89168 99748 89220 99754
rect 89220 99708 89300 99736
rect 89168 99690 89220 99696
rect 88708 99476 88760 99482
rect 88708 99418 88760 99424
rect 88616 98524 88668 98530
rect 88616 98466 88668 98472
rect 88536 98348 88656 98376
rect 88444 97702 88564 97730
rect 88432 97640 88484 97646
rect 88432 97582 88484 97588
rect 88340 94580 88392 94586
rect 88340 94522 88392 94528
rect 88340 94444 88392 94450
rect 88340 94386 88392 94392
rect 88168 16546 88288 16574
rect 87800 6886 88012 6914
rect 87696 4820 87748 4826
rect 87696 4762 87748 4768
rect 87604 4004 87656 4010
rect 87604 3946 87656 3952
rect 87420 3460 87472 3466
rect 87420 3402 87472 3408
rect 87144 3188 87196 3194
rect 87144 3130 87196 3136
rect 87800 490 87828 6886
rect 81594 326 81848 354
rect 81594 -960 81706 326
rect 82698 -960 82810 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86010 -960 86122 480
rect 87114 354 87226 480
rect 87616 462 87828 490
rect 88260 480 88288 16546
rect 88352 3874 88380 94386
rect 88444 4146 88472 97582
rect 88536 94500 88564 97702
rect 88628 94602 88656 98348
rect 88720 94790 88748 99418
rect 88708 94784 88760 94790
rect 88708 94726 88760 94732
rect 88812 94722 88840 99606
rect 88892 98524 88944 98530
rect 88892 98466 88944 98472
rect 88800 94716 88852 94722
rect 88800 94658 88852 94664
rect 88628 94574 88840 94602
rect 88536 94472 88748 94500
rect 88524 94376 88576 94382
rect 88524 94318 88576 94324
rect 88616 94376 88668 94382
rect 88616 94318 88668 94324
rect 88432 4140 88484 4146
rect 88432 4082 88484 4088
rect 88340 3868 88392 3874
rect 88340 3810 88392 3816
rect 88536 3398 88564 94318
rect 88628 3738 88656 94318
rect 88720 4350 88748 94472
rect 88708 4344 88760 4350
rect 88708 4286 88760 4292
rect 88812 4214 88840 94574
rect 88904 5302 88932 98466
rect 88996 5506 89024 99622
rect 89088 99606 89208 99634
rect 89076 99544 89128 99550
rect 89076 99486 89128 99492
rect 89088 97646 89116 99486
rect 89076 97640 89128 97646
rect 89076 97582 89128 97588
rect 89076 94784 89128 94790
rect 89076 94726 89128 94732
rect 89088 19990 89116 94726
rect 89180 46306 89208 99606
rect 89272 98394 89300 99708
rect 89364 99657 89392 99776
rect 89686 99804 89714 100028
rect 89490 99758 89542 99764
rect 89640 99776 89714 99804
rect 89444 99680 89496 99686
rect 89350 99648 89406 99657
rect 89444 99622 89496 99628
rect 89536 99680 89588 99686
rect 89536 99622 89588 99628
rect 89350 99583 89406 99592
rect 89352 99408 89404 99414
rect 89352 99350 89404 99356
rect 89260 98388 89312 98394
rect 89260 98330 89312 98336
rect 89168 46300 89220 46306
rect 89168 46242 89220 46248
rect 89076 19984 89128 19990
rect 89076 19926 89128 19932
rect 88984 5500 89036 5506
rect 88984 5442 89036 5448
rect 88892 5296 88944 5302
rect 88892 5238 88944 5244
rect 88800 4208 88852 4214
rect 88800 4150 88852 4156
rect 88616 3732 88668 3738
rect 88616 3674 88668 3680
rect 89364 3534 89392 99350
rect 89456 98190 89484 99622
rect 89444 98184 89496 98190
rect 89444 98126 89496 98132
rect 89548 97170 89576 99622
rect 89640 98025 89668 99776
rect 89778 99736 89806 100028
rect 89870 99963 89898 100028
rect 89856 99954 89912 99963
rect 89856 99889 89912 99898
rect 89732 99708 89806 99736
rect 89732 98326 89760 99708
rect 89962 99668 89990 100028
rect 90054 99929 90082 100028
rect 90040 99920 90096 99929
rect 90040 99855 90096 99864
rect 90146 99668 90174 100028
rect 90238 99890 90266 100028
rect 90330 99958 90358 100028
rect 90422 99958 90450 100028
rect 90606 99958 90634 100028
rect 90318 99952 90370 99958
rect 90318 99894 90370 99900
rect 90410 99952 90462 99958
rect 90410 99894 90462 99900
rect 90594 99952 90646 99958
rect 90698 99929 90726 100028
rect 90594 99894 90646 99900
rect 90684 99920 90740 99929
rect 90226 99884 90278 99890
rect 90684 99855 90740 99864
rect 90226 99826 90278 99832
rect 90640 99816 90692 99822
rect 90790 99793 90818 100028
rect 90640 99758 90692 99764
rect 90776 99784 90832 99793
rect 90364 99748 90416 99754
rect 89810 99648 89866 99657
rect 89962 99640 90036 99668
rect 89810 99583 89866 99592
rect 89720 98320 89772 98326
rect 89720 98262 89772 98268
rect 89720 98184 89772 98190
rect 89720 98126 89772 98132
rect 89626 98016 89682 98025
rect 89626 97951 89682 97960
rect 89626 97880 89682 97889
rect 89626 97815 89682 97824
rect 89536 97164 89588 97170
rect 89536 97106 89588 97112
rect 89640 94382 89668 97815
rect 89628 94376 89680 94382
rect 89628 94318 89680 94324
rect 89732 5234 89760 98126
rect 89824 94450 89852 99583
rect 89904 99544 89956 99550
rect 89904 99486 89956 99492
rect 89916 98433 89944 99486
rect 89902 98424 89958 98433
rect 89902 98359 89958 98368
rect 89904 98320 89956 98326
rect 89904 98262 89956 98268
rect 89916 94602 89944 98262
rect 90008 97714 90036 99640
rect 90100 99640 90174 99668
rect 90284 99708 90364 99736
rect 90100 98122 90128 99640
rect 90178 98288 90234 98297
rect 90178 98223 90234 98232
rect 90088 98116 90140 98122
rect 90088 98058 90140 98064
rect 89996 97708 90048 97714
rect 89996 97650 90048 97656
rect 89916 94574 90036 94602
rect 89904 94512 89956 94518
rect 89904 94454 89956 94460
rect 89812 94444 89864 94450
rect 89812 94386 89864 94392
rect 89812 94308 89864 94314
rect 89812 94250 89864 94256
rect 89720 5228 89772 5234
rect 89720 5170 89772 5176
rect 89352 3528 89404 3534
rect 89352 3470 89404 3476
rect 88524 3392 88576 3398
rect 88524 3334 88576 3340
rect 89824 3330 89852 94250
rect 89916 4826 89944 94454
rect 90008 5098 90036 94574
rect 90088 94580 90140 94586
rect 90088 94522 90140 94528
rect 90100 6186 90128 94522
rect 90192 6254 90220 98223
rect 90284 94586 90312 99708
rect 90364 99690 90416 99696
rect 90548 99680 90600 99686
rect 90362 99648 90418 99657
rect 90548 99622 90600 99628
rect 90362 99583 90418 99592
rect 90272 94580 90324 94586
rect 90272 94522 90324 94528
rect 90272 94444 90324 94450
rect 90272 94386 90324 94392
rect 90284 21418 90312 94386
rect 90376 91798 90404 99583
rect 90456 97164 90508 97170
rect 90456 97106 90508 97112
rect 90364 91792 90416 91798
rect 90364 91734 90416 91740
rect 90272 21412 90324 21418
rect 90272 21354 90324 21360
rect 90180 6248 90232 6254
rect 90180 6190 90232 6196
rect 90088 6180 90140 6186
rect 90088 6122 90140 6128
rect 90468 5166 90496 97106
rect 90560 94314 90588 99622
rect 90652 94518 90680 99758
rect 90776 99719 90832 99728
rect 90730 99648 90786 99657
rect 90882 99634 90910 100028
rect 90974 99963 91002 100028
rect 90960 99954 91016 99963
rect 90960 99889 91016 99898
rect 91066 99736 91094 100028
rect 91158 99804 91186 100028
rect 91250 99958 91278 100028
rect 91238 99952 91290 99958
rect 91238 99894 91290 99900
rect 91342 99822 91370 100028
rect 91330 99816 91382 99822
rect 91158 99793 91232 99804
rect 91158 99784 91246 99793
rect 91158 99776 91190 99784
rect 91066 99708 91140 99736
rect 91330 99758 91382 99764
rect 91190 99719 91246 99728
rect 91434 99736 91462 100028
rect 91526 99890 91554 100028
rect 91618 99890 91646 100028
rect 91514 99884 91566 99890
rect 91514 99826 91566 99832
rect 91606 99884 91658 99890
rect 91606 99826 91658 99832
rect 91710 99736 91738 100028
rect 91802 99958 91830 100028
rect 91894 99963 91922 100028
rect 91790 99952 91842 99958
rect 91790 99894 91842 99900
rect 91880 99954 91936 99963
rect 91880 99889 91936 99898
rect 91834 99784 91890 99793
rect 91434 99708 91508 99736
rect 91710 99708 91784 99736
rect 91986 99736 92014 100028
rect 91834 99719 91890 99728
rect 90786 99606 90910 99634
rect 91008 99612 91060 99618
rect 90730 99583 90786 99592
rect 91008 99554 91060 99560
rect 90732 99476 90784 99482
rect 90732 99418 90784 99424
rect 90640 94512 90692 94518
rect 90640 94454 90692 94460
rect 90548 94308 90600 94314
rect 90548 94250 90600 94256
rect 90456 5160 90508 5166
rect 90456 5102 90508 5108
rect 89996 5092 90048 5098
rect 89996 5034 90048 5040
rect 89904 4820 89956 4826
rect 89904 4762 89956 4768
rect 90744 3602 90772 99418
rect 90824 99408 90876 99414
rect 90824 99350 90876 99356
rect 90836 97442 90864 99350
rect 90916 98388 90968 98394
rect 90916 98330 90968 98336
rect 90824 97436 90876 97442
rect 90824 97378 90876 97384
rect 90928 84194 90956 98330
rect 91020 97238 91048 99554
rect 91112 97918 91140 99708
rect 91192 99680 91244 99686
rect 91192 99622 91244 99628
rect 91374 99648 91430 99657
rect 91100 97912 91152 97918
rect 91100 97854 91152 97860
rect 91100 97708 91152 97714
rect 91100 97650 91152 97656
rect 91008 97232 91060 97238
rect 91008 97174 91060 97180
rect 91112 94450 91140 97650
rect 91100 94444 91152 94450
rect 91100 94386 91152 94392
rect 90836 84166 90956 84194
rect 90836 5370 90864 84166
rect 91204 6594 91232 99622
rect 91284 99612 91336 99618
rect 91374 99583 91430 99592
rect 91284 99554 91336 99560
rect 91296 94994 91324 99554
rect 91388 95234 91416 99583
rect 91480 98190 91508 99708
rect 91652 99612 91704 99618
rect 91572 99572 91652 99600
rect 91468 98184 91520 98190
rect 91468 98126 91520 98132
rect 91572 97102 91600 99572
rect 91652 99554 91704 99560
rect 91756 98240 91784 99708
rect 91664 98212 91784 98240
rect 91664 97714 91692 98212
rect 91744 98116 91796 98122
rect 91744 98058 91796 98064
rect 91652 97708 91704 97714
rect 91652 97650 91704 97656
rect 91560 97096 91612 97102
rect 91560 97038 91612 97044
rect 91388 95206 91508 95234
rect 91284 94988 91336 94994
rect 91284 94930 91336 94936
rect 91376 94648 91428 94654
rect 91376 94590 91428 94596
rect 91284 94580 91336 94586
rect 91284 94522 91336 94528
rect 91296 42090 91324 94522
rect 91388 87650 91416 94590
rect 91480 90370 91508 95206
rect 91468 90364 91520 90370
rect 91468 90306 91520 90312
rect 91376 87644 91428 87650
rect 91376 87586 91428 87592
rect 91284 42084 91336 42090
rect 91284 42026 91336 42032
rect 91192 6588 91244 6594
rect 91192 6530 91244 6536
rect 91756 6322 91784 98058
rect 91848 94654 91876 99719
rect 91940 99708 92014 99736
rect 92078 99736 92106 100028
rect 92170 99890 92198 100028
rect 92262 99963 92290 100028
rect 92248 99954 92304 99963
rect 92354 99958 92382 100028
rect 92158 99884 92210 99890
rect 92248 99889 92304 99898
rect 92342 99952 92394 99958
rect 92342 99894 92394 99900
rect 92446 99890 92474 100028
rect 92158 99826 92210 99832
rect 92434 99884 92486 99890
rect 92434 99826 92486 99832
rect 92538 99736 92566 100028
rect 92630 99963 92658 100028
rect 92616 99954 92672 99963
rect 92722 99958 92750 100028
rect 92616 99889 92672 99898
rect 92710 99952 92762 99958
rect 92710 99894 92762 99900
rect 92814 99895 92842 100028
rect 92906 99958 92934 100028
rect 92998 99958 93026 100028
rect 92894 99952 92946 99958
rect 92800 99886 92856 99895
rect 92894 99894 92946 99900
rect 92986 99952 93038 99958
rect 92986 99894 93038 99900
rect 92800 99821 92856 99830
rect 93090 99804 93118 100028
rect 92952 99776 93118 99804
rect 92848 99748 92900 99754
rect 92078 99708 92152 99736
rect 92538 99708 92704 99736
rect 91836 94648 91888 94654
rect 91836 94590 91888 94596
rect 91940 94586 91968 99708
rect 92020 99612 92072 99618
rect 92020 99554 92072 99560
rect 92032 97782 92060 99554
rect 92124 98002 92152 99708
rect 92296 99680 92348 99686
rect 92216 99628 92296 99634
rect 92216 99622 92348 99628
rect 92570 99648 92626 99657
rect 92216 99606 92336 99622
rect 92480 99612 92532 99618
rect 92216 98161 92244 99606
rect 92570 99583 92626 99592
rect 92480 99554 92532 99560
rect 92296 99544 92348 99550
rect 92348 99504 92428 99532
rect 92296 99486 92348 99492
rect 92202 98152 92258 98161
rect 92202 98087 92258 98096
rect 92294 98016 92350 98025
rect 92124 97974 92244 98002
rect 92112 97912 92164 97918
rect 92112 97854 92164 97860
rect 92020 97776 92072 97782
rect 92020 97718 92072 97724
rect 92020 97436 92072 97442
rect 92020 97378 92072 97384
rect 91928 94580 91980 94586
rect 91928 94522 91980 94528
rect 91836 94512 91888 94518
rect 91836 94454 91888 94460
rect 91848 6390 91876 94454
rect 91928 94444 91980 94450
rect 91928 94386 91980 94392
rect 91836 6384 91888 6390
rect 91836 6326 91888 6332
rect 91744 6316 91796 6322
rect 91744 6258 91796 6264
rect 90824 5364 90876 5370
rect 90824 5306 90876 5312
rect 91940 3602 91968 94386
rect 92032 4894 92060 97378
rect 92020 4888 92072 4894
rect 92020 4830 92072 4836
rect 92124 3670 92152 97854
rect 92216 97646 92244 97974
rect 92294 97951 92350 97960
rect 92204 97640 92256 97646
rect 92204 97582 92256 97588
rect 92308 3806 92336 97951
rect 92400 97918 92428 99504
rect 92388 97912 92440 97918
rect 92388 97854 92440 97860
rect 92388 97776 92440 97782
rect 92388 97718 92440 97724
rect 92400 94518 92428 97718
rect 92492 97578 92520 99554
rect 92480 97572 92532 97578
rect 92480 97514 92532 97520
rect 92492 96694 92520 97514
rect 92480 96688 92532 96694
rect 92480 96630 92532 96636
rect 92388 94512 92440 94518
rect 92388 94454 92440 94460
rect 92584 94382 92612 99583
rect 92572 94376 92624 94382
rect 92572 94318 92624 94324
rect 92572 94240 92624 94246
rect 92572 94182 92624 94188
rect 92584 89622 92612 94182
rect 92572 89616 92624 89622
rect 92572 89558 92624 89564
rect 92676 24546 92704 99708
rect 92848 99690 92900 99696
rect 92754 99648 92810 99657
rect 92754 99583 92810 99592
rect 92768 26110 92796 99583
rect 92860 97578 92888 99690
rect 92848 97572 92900 97578
rect 92848 97514 92900 97520
rect 92952 94602 92980 99776
rect 93182 99736 93210 100028
rect 93274 99958 93302 100028
rect 93366 99958 93394 100028
rect 93262 99952 93314 99958
rect 93262 99894 93314 99900
rect 93354 99952 93406 99958
rect 93354 99894 93406 99900
rect 93308 99816 93360 99822
rect 93458 99793 93486 100028
rect 93308 99758 93360 99764
rect 93444 99784 93500 99793
rect 92860 94574 92980 94602
rect 93044 99708 93210 99736
rect 92860 27334 92888 94574
rect 93044 94466 93072 99708
rect 93320 99657 93348 99758
rect 93444 99719 93500 99728
rect 93550 99736 93578 100028
rect 93642 99963 93670 100028
rect 93628 99954 93684 99963
rect 93826 99940 93854 100028
rect 93918 99958 93946 100028
rect 94010 99958 94038 100028
rect 93628 99889 93684 99898
rect 93780 99912 93854 99940
rect 93906 99952 93958 99958
rect 93550 99708 93624 99736
rect 93400 99680 93452 99686
rect 93306 99648 93362 99657
rect 93124 99612 93176 99618
rect 93124 99554 93176 99560
rect 93216 99612 93268 99618
rect 93400 99622 93452 99628
rect 93306 99583 93362 99592
rect 93216 99554 93268 99560
rect 93136 97617 93164 99554
rect 93122 97608 93178 97617
rect 93122 97543 93178 97552
rect 92952 94438 93072 94466
rect 92848 27328 92900 27334
rect 92848 27270 92900 27276
rect 92952 27266 92980 94438
rect 93032 94376 93084 94382
rect 93032 94318 93084 94324
rect 92940 27260 92992 27266
rect 92940 27202 92992 27208
rect 92756 26104 92808 26110
rect 92756 26046 92808 26052
rect 92664 24540 92716 24546
rect 92664 24482 92716 24488
rect 93044 17678 93072 94318
rect 93032 17672 93084 17678
rect 93032 17614 93084 17620
rect 93136 10810 93164 97543
rect 93228 96082 93256 99554
rect 93308 99476 93360 99482
rect 93308 99418 93360 99424
rect 93216 96076 93268 96082
rect 93216 96018 93268 96024
rect 93228 12238 93256 96018
rect 93320 95878 93348 99418
rect 93412 98297 93440 99622
rect 93596 99482 93624 99708
rect 93674 99648 93730 99657
rect 93674 99583 93730 99592
rect 93584 99476 93636 99482
rect 93584 99418 93636 99424
rect 93584 99340 93636 99346
rect 93584 99282 93636 99288
rect 93398 98288 93454 98297
rect 93398 98223 93454 98232
rect 93596 97714 93624 99282
rect 93584 97708 93636 97714
rect 93584 97650 93636 97656
rect 93688 97594 93716 99583
rect 93492 97572 93544 97578
rect 93492 97514 93544 97520
rect 93596 97566 93716 97594
rect 93400 97300 93452 97306
rect 93400 97242 93452 97248
rect 93412 96830 93440 97242
rect 93400 96824 93452 96830
rect 93400 96766 93452 96772
rect 93400 96688 93452 96694
rect 93400 96630 93452 96636
rect 93308 95872 93360 95878
rect 93308 95814 93360 95820
rect 93320 13530 93348 95814
rect 93412 92410 93440 96630
rect 93400 92404 93452 92410
rect 93400 92346 93452 92352
rect 93504 89714 93532 97514
rect 93596 95810 93624 97566
rect 93676 97232 93728 97238
rect 93676 97174 93728 97180
rect 93584 95804 93636 95810
rect 93584 95746 93636 95752
rect 93688 94246 93716 97174
rect 93780 96354 93808 99912
rect 93906 99894 93958 99900
rect 93998 99952 94050 99958
rect 93998 99894 94050 99900
rect 94102 99736 94130 100028
rect 94056 99708 94130 99736
rect 93860 99680 93912 99686
rect 94056 99657 94084 99708
rect 94194 99668 94222 100028
rect 94286 99736 94314 100028
rect 94378 99958 94406 100028
rect 94366 99952 94418 99958
rect 94366 99894 94418 99900
rect 94470 99804 94498 100028
rect 94562 99890 94590 100028
rect 94654 99958 94682 100028
rect 94746 99958 94774 100028
rect 94642 99952 94694 99958
rect 94642 99894 94694 99900
rect 94734 99952 94786 99958
rect 94838 99929 94866 100028
rect 94930 99958 94958 100028
rect 94918 99952 94970 99958
rect 94734 99894 94786 99900
rect 94824 99920 94880 99929
rect 94550 99884 94602 99890
rect 94918 99894 94970 99900
rect 94824 99855 94880 99864
rect 94550 99826 94602 99832
rect 94424 99776 94498 99804
rect 94688 99816 94740 99822
rect 94686 99784 94688 99793
rect 95022 99793 95050 100028
rect 95114 99890 95142 100028
rect 95102 99884 95154 99890
rect 95102 99826 95154 99832
rect 95206 99822 95234 100028
rect 95194 99816 95246 99822
rect 94740 99784 94742 99793
rect 94286 99708 94360 99736
rect 93860 99622 93912 99628
rect 94042 99648 94098 99657
rect 93768 96348 93820 96354
rect 93768 96290 93820 96296
rect 93872 94738 93900 99622
rect 93952 99612 94004 99618
rect 94042 99583 94098 99592
rect 94148 99640 94222 99668
rect 93952 99554 94004 99560
rect 93780 94710 93900 94738
rect 93780 94450 93808 94710
rect 93860 94580 93912 94586
rect 93860 94522 93912 94528
rect 93768 94444 93820 94450
rect 93768 94386 93820 94392
rect 93676 94240 93728 94246
rect 93676 94182 93728 94188
rect 93504 89686 93624 89714
rect 93596 21894 93624 89686
rect 93584 21888 93636 21894
rect 93584 21830 93636 21836
rect 93872 18970 93900 94522
rect 93964 30190 93992 99554
rect 94044 99544 94096 99550
rect 94044 99486 94096 99492
rect 94056 94586 94084 99486
rect 94044 94580 94096 94586
rect 94044 94522 94096 94528
rect 94044 94444 94096 94450
rect 94044 94386 94096 94392
rect 94056 31550 94084 94386
rect 94044 31544 94096 31550
rect 94044 31486 94096 31492
rect 94148 31482 94176 99640
rect 94228 99544 94280 99550
rect 94228 99486 94280 99492
rect 94240 96422 94268 99486
rect 94228 96416 94280 96422
rect 94228 96358 94280 96364
rect 94228 94580 94280 94586
rect 94228 94522 94280 94528
rect 94240 41206 94268 94522
rect 94332 85202 94360 99708
rect 94424 94586 94452 99776
rect 95008 99784 95064 99793
rect 94686 99719 94742 99728
rect 94872 99748 94924 99754
rect 95194 99758 95246 99764
rect 95008 99719 95064 99728
rect 94872 99690 94924 99696
rect 94780 97096 94832 97102
rect 94780 97038 94832 97044
rect 94688 96416 94740 96422
rect 94688 96358 94740 96364
rect 94596 96348 94648 96354
rect 94596 96290 94648 96296
rect 94504 95804 94556 95810
rect 94504 95746 94556 95752
rect 94412 94580 94464 94586
rect 94412 94522 94464 94528
rect 94516 89714 94544 95746
rect 94608 90710 94636 96290
rect 94596 90704 94648 90710
rect 94596 90646 94648 90652
rect 94516 89686 94636 89714
rect 94502 88224 94558 88233
rect 94502 88159 94558 88168
rect 94320 85196 94372 85202
rect 94320 85138 94372 85144
rect 94228 41200 94280 41206
rect 94228 41142 94280 41148
rect 94136 31476 94188 31482
rect 94136 31418 94188 31424
rect 93952 30184 94004 30190
rect 93952 30126 94004 30132
rect 93860 18964 93912 18970
rect 93860 18906 93912 18912
rect 93308 13524 93360 13530
rect 93308 13466 93360 13472
rect 93216 12232 93268 12238
rect 93216 12174 93268 12180
rect 93124 10804 93176 10810
rect 93124 10746 93176 10752
rect 93768 4208 93820 4214
rect 93768 4150 93820 4156
rect 92296 3800 92348 3806
rect 92296 3742 92348 3748
rect 92112 3664 92164 3670
rect 92112 3606 92164 3612
rect 90732 3596 90784 3602
rect 90732 3538 90784 3544
rect 91928 3596 91980 3602
rect 91928 3538 91980 3544
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 90456 3460 90508 3466
rect 90456 3402 90508 3408
rect 89812 3324 89864 3330
rect 89812 3266 89864 3272
rect 89352 3188 89404 3194
rect 89352 3130 89404 3136
rect 89364 480 89392 3130
rect 90468 480 90496 3402
rect 91572 480 91600 3470
rect 92664 3392 92716 3398
rect 92664 3334 92716 3340
rect 92676 480 92704 3334
rect 93780 480 93808 4150
rect 94516 3942 94544 88159
rect 94608 16318 94636 89686
rect 94700 17610 94728 96358
rect 94792 42158 94820 97038
rect 94884 96490 94912 99690
rect 94964 99680 95016 99686
rect 95298 99668 95326 100028
rect 95390 99804 95418 100028
rect 95482 99929 95510 100028
rect 95468 99920 95524 99929
rect 95468 99855 95524 99864
rect 95574 99804 95602 100028
rect 95666 99963 95694 100028
rect 95652 99954 95708 99963
rect 95758 99958 95786 100028
rect 95652 99889 95708 99898
rect 95746 99952 95798 99958
rect 95746 99894 95798 99900
rect 95390 99776 95464 99804
rect 94964 99622 95016 99628
rect 95252 99640 95326 99668
rect 94976 97238 95004 99622
rect 95056 99476 95108 99482
rect 95056 99418 95108 99424
rect 95148 99476 95200 99482
rect 95148 99418 95200 99424
rect 95068 97306 95096 99418
rect 95160 97889 95188 99418
rect 95252 98530 95280 99640
rect 95436 99464 95464 99776
rect 95528 99776 95602 99804
rect 95652 99784 95708 99793
rect 95528 99668 95556 99776
rect 95850 99770 95878 100028
rect 95942 99958 95970 100028
rect 96034 99958 96062 100028
rect 95930 99952 95982 99958
rect 95930 99894 95982 99900
rect 96022 99952 96074 99958
rect 96022 99894 96074 99900
rect 95804 99742 95878 99770
rect 95976 99816 96028 99822
rect 95976 99758 96028 99764
rect 95708 99728 95740 99736
rect 95652 99719 95740 99728
rect 95666 99708 95740 99719
rect 95528 99640 95648 99668
rect 95344 99436 95464 99464
rect 95240 98524 95292 98530
rect 95240 98466 95292 98472
rect 95344 98376 95372 99436
rect 95424 98524 95476 98530
rect 95424 98466 95476 98472
rect 95252 98348 95372 98376
rect 95146 97880 95202 97889
rect 95146 97815 95202 97824
rect 95056 97300 95108 97306
rect 95056 97242 95108 97248
rect 94964 97232 95016 97238
rect 94964 97174 95016 97180
rect 94872 96484 94924 96490
rect 94872 96426 94924 96432
rect 95252 96354 95280 98348
rect 95330 98288 95386 98297
rect 95330 98223 95386 98232
rect 95344 96626 95372 98223
rect 95332 96620 95384 96626
rect 95332 96562 95384 96568
rect 95240 96348 95292 96354
rect 95240 96290 95292 96296
rect 95344 95266 95372 96562
rect 95332 95260 95384 95266
rect 95332 95202 95384 95208
rect 94780 42152 94832 42158
rect 94780 42094 94832 42100
rect 95436 21826 95464 98466
rect 95516 94580 95568 94586
rect 95516 94522 95568 94528
rect 95528 23118 95556 94522
rect 95620 23186 95648 99640
rect 95712 36718 95740 99708
rect 95804 94586 95832 99742
rect 95884 99680 95936 99686
rect 95884 99622 95936 99628
rect 95896 94722 95924 99622
rect 95988 96218 96016 99758
rect 96126 99736 96154 100028
rect 96218 99929 96246 100028
rect 96310 99958 96338 100028
rect 96298 99952 96350 99958
rect 96204 99920 96260 99929
rect 96298 99894 96350 99900
rect 96204 99855 96260 99864
rect 96402 99793 96430 100028
rect 96388 99784 96444 99793
rect 96126 99708 96292 99736
rect 96388 99719 96444 99728
rect 96068 99272 96120 99278
rect 96068 99214 96120 99220
rect 95976 96212 96028 96218
rect 95976 96154 96028 96160
rect 95884 94716 95936 94722
rect 95884 94658 95936 94664
rect 95792 94580 95844 94586
rect 95792 94522 95844 94528
rect 95884 94580 95936 94586
rect 95884 94522 95936 94528
rect 95896 89486 95924 94522
rect 95988 94466 96016 96154
rect 96080 94586 96108 99214
rect 96160 95260 96212 95266
rect 96160 95202 96212 95208
rect 96068 94580 96120 94586
rect 96068 94522 96120 94528
rect 95988 94438 96108 94466
rect 95976 94376 96028 94382
rect 95976 94318 96028 94324
rect 95884 89480 95936 89486
rect 95884 89422 95936 89428
rect 95700 36712 95752 36718
rect 95700 36654 95752 36660
rect 95608 23180 95660 23186
rect 95608 23122 95660 23128
rect 95516 23112 95568 23118
rect 95516 23054 95568 23060
rect 95424 21820 95476 21826
rect 95424 21762 95476 21768
rect 94688 17604 94740 17610
rect 94688 17546 94740 17552
rect 94596 16312 94648 16318
rect 94596 16254 94648 16260
rect 95988 6458 96016 94318
rect 96080 6526 96108 94438
rect 96172 89554 96200 95202
rect 96160 89548 96212 89554
rect 96160 89490 96212 89496
rect 96068 6520 96120 6526
rect 96068 6462 96120 6468
rect 95976 6452 96028 6458
rect 95976 6394 96028 6400
rect 96264 5438 96292 99708
rect 96494 99668 96522 100028
rect 96586 99958 96614 100028
rect 96574 99952 96626 99958
rect 96574 99894 96626 99900
rect 96678 99804 96706 100028
rect 96770 99929 96798 100028
rect 96756 99920 96812 99929
rect 96862 99890 96890 100028
rect 96954 99958 96982 100028
rect 97046 99963 97074 100028
rect 96942 99952 96994 99958
rect 96942 99894 96994 99900
rect 97032 99954 97088 99963
rect 96756 99855 96812 99864
rect 96850 99884 96902 99890
rect 97032 99889 97088 99898
rect 97138 99890 97166 100028
rect 97230 99963 97258 100028
rect 97216 99954 97272 99963
rect 96850 99826 96902 99832
rect 97126 99884 97178 99890
rect 97216 99889 97272 99898
rect 97322 99890 97350 100028
rect 97414 99963 97442 100028
rect 97400 99954 97456 99963
rect 97506 99940 97534 100028
rect 97690 99958 97718 100028
rect 97678 99952 97730 99958
rect 97506 99912 97580 99940
rect 97126 99826 97178 99832
rect 97310 99884 97362 99890
rect 97400 99889 97456 99898
rect 97310 99826 97362 99832
rect 96678 99776 96798 99804
rect 97552 99793 97580 99912
rect 97678 99894 97730 99900
rect 97782 99890 97810 100028
rect 97770 99884 97822 99890
rect 97770 99826 97822 99832
rect 96770 99770 96798 99776
rect 97354 99784 97410 99793
rect 96770 99742 96844 99770
rect 96712 99680 96764 99686
rect 96494 99640 96568 99668
rect 96436 99544 96488 99550
rect 96436 99486 96488 99492
rect 96448 96286 96476 99486
rect 96540 97617 96568 99640
rect 96618 99648 96674 99657
rect 96712 99622 96764 99628
rect 96618 99583 96674 99592
rect 96526 97608 96582 97617
rect 96526 97543 96582 97552
rect 96632 96286 96660 99583
rect 96436 96280 96488 96286
rect 96436 96222 96488 96228
rect 96620 96280 96672 96286
rect 96620 96222 96672 96228
rect 96448 95234 96476 96222
rect 96724 95878 96752 99622
rect 96712 95872 96764 95878
rect 96712 95814 96764 95820
rect 96448 95206 96568 95234
rect 96344 94716 96396 94722
rect 96344 94658 96396 94664
rect 96356 18902 96384 94658
rect 96540 94382 96568 95206
rect 96620 94852 96672 94858
rect 96620 94794 96672 94800
rect 96528 94376 96580 94382
rect 96528 94318 96580 94324
rect 96344 18896 96396 18902
rect 96344 18838 96396 18844
rect 96632 8090 96660 94794
rect 96816 94722 96844 99742
rect 96896 99748 96948 99754
rect 96896 99690 96948 99696
rect 97080 99748 97132 99754
rect 97080 99690 97132 99696
rect 97276 99742 97354 99770
rect 96804 94716 96856 94722
rect 96804 94658 96856 94664
rect 96908 94602 96936 99690
rect 96986 99648 97042 99657
rect 96986 99583 97042 99592
rect 96724 94574 96936 94602
rect 96724 22982 96752 94574
rect 96804 94512 96856 94518
rect 96804 94454 96856 94460
rect 96896 94512 96948 94518
rect 96896 94454 96948 94460
rect 96816 23050 96844 94454
rect 96908 24478 96936 94454
rect 97000 36650 97028 99583
rect 97092 85542 97120 99690
rect 97172 99680 97224 99686
rect 97172 99622 97224 99628
rect 97184 96614 97212 99622
rect 97276 97170 97304 99742
rect 97354 99719 97410 99728
rect 97538 99784 97594 99793
rect 97874 99736 97902 100028
rect 97966 99958 97994 100028
rect 98058 99963 98086 100028
rect 97954 99952 98006 99958
rect 97954 99894 98006 99900
rect 98044 99954 98100 99963
rect 98044 99889 98100 99898
rect 98150 99822 98178 100028
rect 98242 99958 98270 100028
rect 98334 99963 98362 100028
rect 98230 99952 98282 99958
rect 98230 99894 98282 99900
rect 98320 99954 98376 99963
rect 98426 99958 98454 100028
rect 98518 99963 98546 100028
rect 98320 99889 98376 99898
rect 98414 99952 98466 99958
rect 98414 99894 98466 99900
rect 98504 99954 98560 99963
rect 98504 99889 98560 99898
rect 98138 99816 98190 99822
rect 98610 99770 98638 100028
rect 98702 99958 98730 100028
rect 98690 99952 98742 99958
rect 98794 99929 98822 100028
rect 98886 99958 98914 100028
rect 98874 99952 98926 99958
rect 98690 99894 98742 99900
rect 98780 99920 98836 99929
rect 99070 99906 99098 100028
rect 99162 99958 99190 100028
rect 98874 99894 98926 99900
rect 99024 99890 99098 99906
rect 99150 99952 99202 99958
rect 99150 99894 99202 99900
rect 99254 99890 99282 100028
rect 98780 99855 98836 99864
rect 99012 99884 99098 99890
rect 99064 99878 99098 99884
rect 99242 99884 99294 99890
rect 99012 99826 99064 99832
rect 99242 99826 99294 99832
rect 98138 99758 98190 99764
rect 97538 99719 97594 99728
rect 97828 99708 97902 99736
rect 98368 99748 98420 99754
rect 97632 99680 97684 99686
rect 97354 99648 97410 99657
rect 97632 99622 97684 99628
rect 97354 99583 97410 99592
rect 97448 99612 97500 99618
rect 97264 97164 97316 97170
rect 97264 97106 97316 97112
rect 97184 96586 97304 96614
rect 97172 95872 97224 95878
rect 97172 95814 97224 95820
rect 97184 92206 97212 95814
rect 97276 92478 97304 96586
rect 97368 94518 97396 99583
rect 97448 99554 97500 99560
rect 97540 99612 97592 99618
rect 97540 99554 97592 99560
rect 97460 96218 97488 99554
rect 97552 97617 97580 99554
rect 97538 97608 97594 97617
rect 97538 97543 97594 97552
rect 97644 97481 97672 99622
rect 97630 97472 97686 97481
rect 97630 97407 97686 97416
rect 97828 97209 97856 99708
rect 98368 99690 98420 99696
rect 98564 99742 98638 99770
rect 99104 99816 99156 99822
rect 99104 99758 99156 99764
rect 99194 99784 99250 99793
rect 98736 99748 98788 99754
rect 98274 99648 98330 99657
rect 98000 99612 98052 99618
rect 98274 99583 98330 99592
rect 98000 99554 98052 99560
rect 97908 99544 97960 99550
rect 97906 99512 97908 99521
rect 97960 99512 97962 99521
rect 97906 99447 97962 99456
rect 97814 97200 97870 97209
rect 97540 97164 97592 97170
rect 97814 97135 97870 97144
rect 97540 97106 97592 97112
rect 97552 96393 97580 97106
rect 97538 96384 97594 96393
rect 97538 96319 97594 96328
rect 97448 96212 97500 96218
rect 97448 96154 97500 96160
rect 97356 94512 97408 94518
rect 97356 94454 97408 94460
rect 97264 92472 97316 92478
rect 97264 92414 97316 92420
rect 97172 92200 97224 92206
rect 97172 92142 97224 92148
rect 97080 85536 97132 85542
rect 97080 85478 97132 85484
rect 96988 36644 97040 36650
rect 96988 36586 97040 36592
rect 96896 24472 96948 24478
rect 96896 24414 96948 24420
rect 96804 23044 96856 23050
rect 96804 22986 96856 22992
rect 96712 22976 96764 22982
rect 96712 22918 96764 22924
rect 97552 8158 97580 96319
rect 97920 94858 97948 99447
rect 97908 94852 97960 94858
rect 97908 94794 97960 94800
rect 98012 94738 98040 99554
rect 98182 97608 98238 97617
rect 98182 97543 98238 97552
rect 98090 97064 98146 97073
rect 98090 96999 98146 97008
rect 97920 94710 98040 94738
rect 98104 94722 98132 96999
rect 98092 94716 98144 94722
rect 97920 94314 97948 94710
rect 98092 94658 98144 94664
rect 98000 94648 98052 94654
rect 98000 94590 98052 94596
rect 97908 94308 97960 94314
rect 97908 94250 97960 94256
rect 98012 20466 98040 94590
rect 98092 94580 98144 94586
rect 98092 94522 98144 94528
rect 98104 24342 98132 94522
rect 98196 24410 98224 97543
rect 98288 94586 98316 99583
rect 98380 94654 98408 99690
rect 98460 99680 98512 99686
rect 98460 99622 98512 99628
rect 98472 97850 98500 99622
rect 98460 97844 98512 97850
rect 98460 97786 98512 97792
rect 98564 97730 98592 99742
rect 98736 99690 98788 99696
rect 98920 99748 98972 99754
rect 98920 99690 98972 99696
rect 98642 99648 98698 99657
rect 98642 99583 98698 99592
rect 98656 97753 98684 99583
rect 98472 97702 98592 97730
rect 98642 97744 98698 97753
rect 98368 94648 98420 94654
rect 98368 94590 98420 94596
rect 98276 94580 98328 94586
rect 98276 94522 98328 94528
rect 98472 94466 98500 97702
rect 98642 97679 98698 97688
rect 98552 97572 98604 97578
rect 98552 97514 98604 97520
rect 98288 94438 98500 94466
rect 98184 24404 98236 24410
rect 98184 24346 98236 24352
rect 98092 24336 98144 24342
rect 98092 24278 98144 24284
rect 98288 24274 98316 94438
rect 98368 94376 98420 94382
rect 98368 94318 98420 94324
rect 98380 32910 98408 94318
rect 98460 94308 98512 94314
rect 98460 94250 98512 94256
rect 98472 88330 98500 94250
rect 98564 89690 98592 97514
rect 98656 89714 98684 97679
rect 98748 94382 98776 99690
rect 98828 99612 98880 99618
rect 98828 99554 98880 99560
rect 98840 99521 98868 99554
rect 98826 99512 98882 99521
rect 98826 99447 98882 99456
rect 98828 97844 98880 97850
rect 98828 97786 98880 97792
rect 98736 94376 98788 94382
rect 98736 94318 98788 94324
rect 98840 91050 98868 97786
rect 98932 97617 98960 99690
rect 99012 99476 99064 99482
rect 99012 99418 99064 99424
rect 98918 97608 98974 97617
rect 98918 97543 98974 97552
rect 99024 97481 99052 99418
rect 99116 97617 99144 99758
rect 99194 99719 99250 99728
rect 99346 99736 99374 100028
rect 99438 99890 99466 100028
rect 99530 99958 99558 100028
rect 99518 99952 99570 99958
rect 99714 99929 99742 100028
rect 99518 99894 99570 99900
rect 99700 99920 99756 99929
rect 99426 99884 99478 99890
rect 99700 99855 99756 99864
rect 99426 99826 99478 99832
rect 99656 99816 99708 99822
rect 99654 99784 99656 99793
rect 99708 99784 99710 99793
rect 99564 99748 99616 99754
rect 99102 97608 99158 97617
rect 99208 97578 99236 99719
rect 99346 99708 99512 99736
rect 99286 99648 99342 99657
rect 99286 99583 99342 99592
rect 99102 97543 99158 97552
rect 99196 97572 99248 97578
rect 99196 97514 99248 97520
rect 99010 97472 99066 97481
rect 99010 97407 99066 97416
rect 99300 96614 99328 99583
rect 99300 96586 99420 96614
rect 99288 94716 99340 94722
rect 99288 94658 99340 94664
rect 98828 91044 98880 91050
rect 98828 90986 98880 90992
rect 98552 89684 98604 89690
rect 98656 89686 98960 89714
rect 98552 89626 98604 89632
rect 98642 89040 98698 89049
rect 98642 88975 98698 88984
rect 98460 88324 98512 88330
rect 98460 88266 98512 88272
rect 98368 32904 98420 32910
rect 98368 32846 98420 32852
rect 98276 24268 98328 24274
rect 98276 24210 98328 24216
rect 98000 20460 98052 20466
rect 98000 20402 98052 20408
rect 98092 19984 98144 19990
rect 98092 19926 98144 19932
rect 98104 16574 98132 19926
rect 98104 16546 98224 16574
rect 97540 8152 97592 8158
rect 97540 8094 97592 8100
rect 96620 8084 96672 8090
rect 96620 8026 96672 8032
rect 96252 5432 96304 5438
rect 96252 5374 96304 5380
rect 97080 5296 97132 5302
rect 97080 5238 97132 5244
rect 94872 4344 94924 4350
rect 94872 4286 94924 4292
rect 94504 3936 94556 3942
rect 94504 3878 94556 3884
rect 94884 480 94912 4286
rect 95976 4140 96028 4146
rect 95976 4082 96028 4088
rect 95988 480 96016 4082
rect 97092 480 97120 5238
rect 98196 480 98224 16546
rect 98656 4078 98684 88975
rect 98932 84194 98960 89686
rect 98840 84166 98960 84194
rect 98840 8022 98868 84166
rect 98828 8016 98880 8022
rect 98828 7958 98880 7964
rect 99300 7954 99328 94658
rect 99392 89714 99420 96586
rect 99484 92138 99512 99708
rect 99654 99719 99710 99728
rect 99564 99690 99616 99696
rect 99472 92132 99524 92138
rect 99472 92074 99524 92080
rect 99392 89686 99512 89714
rect 99288 7948 99340 7954
rect 99288 7890 99340 7896
rect 99484 7886 99512 89686
rect 99576 21758 99604 99690
rect 99806 99668 99834 100028
rect 99898 99770 99926 100028
rect 99990 99929 100018 100028
rect 99976 99920 100032 99929
rect 100082 99890 100110 100028
rect 100174 99958 100202 100028
rect 100266 99958 100294 100028
rect 100162 99952 100214 99958
rect 100162 99894 100214 99900
rect 100254 99952 100306 99958
rect 100358 99929 100386 100028
rect 100450 99958 100478 100028
rect 100438 99952 100490 99958
rect 100254 99894 100306 99900
rect 100344 99920 100400 99929
rect 99976 99855 100032 99864
rect 100070 99884 100122 99890
rect 100070 99826 100122 99832
rect 100174 99804 100202 99894
rect 100438 99894 100490 99900
rect 100344 99855 100400 99864
rect 100174 99776 100432 99804
rect 99898 99742 100064 99770
rect 99668 99640 99834 99668
rect 99668 38282 99696 99640
rect 99932 99612 99984 99618
rect 99932 99554 99984 99560
rect 99748 99544 99800 99550
rect 99748 99486 99800 99492
rect 99656 38276 99708 38282
rect 99656 38218 99708 38224
rect 99760 38214 99788 99486
rect 99840 99476 99892 99482
rect 99840 99418 99892 99424
rect 99852 46238 99880 99418
rect 99944 88262 99972 99554
rect 100036 99482 100064 99742
rect 100114 99648 100170 99657
rect 100114 99583 100170 99592
rect 100208 99612 100260 99618
rect 100024 99476 100076 99482
rect 100024 99418 100076 99424
rect 100036 94586 100064 99418
rect 100024 94580 100076 94586
rect 100024 94522 100076 94528
rect 99932 88256 99984 88262
rect 99932 88198 99984 88204
rect 100024 46300 100076 46306
rect 100024 46242 100076 46248
rect 99840 46232 99892 46238
rect 99840 46174 99892 46180
rect 99748 38208 99800 38214
rect 99748 38150 99800 38156
rect 99564 21752 99616 21758
rect 99564 21694 99616 21700
rect 99472 7880 99524 7886
rect 99472 7822 99524 7828
rect 98644 4072 98696 4078
rect 98644 4014 98696 4020
rect 99288 3868 99340 3874
rect 99288 3810 99340 3816
rect 99300 480 99328 3810
rect 100036 3398 100064 46242
rect 100128 5302 100156 99583
rect 100208 99554 100260 99560
rect 100220 98297 100248 99554
rect 100206 98288 100262 98297
rect 100206 98223 100262 98232
rect 100404 96614 100432 99776
rect 100542 99736 100570 100028
rect 100634 99958 100662 100028
rect 100622 99952 100674 99958
rect 100818 99906 100846 100028
rect 100910 99958 100938 100028
rect 101002 99963 101030 100028
rect 100622 99894 100674 99900
rect 100772 99878 100846 99906
rect 100898 99952 100950 99958
rect 100898 99894 100950 99900
rect 100988 99954 101044 99963
rect 101094 99958 101122 100028
rect 100988 99889 101044 99898
rect 101082 99952 101134 99958
rect 101082 99894 101134 99900
rect 100668 99816 100720 99822
rect 100668 99758 100720 99764
rect 100542 99708 100616 99736
rect 100484 99612 100536 99618
rect 100484 99554 100536 99560
rect 100312 96586 100432 96614
rect 100312 82346 100340 96586
rect 100496 95234 100524 99554
rect 100588 98161 100616 99708
rect 100680 98433 100708 99758
rect 100772 99634 100800 99878
rect 101186 99770 101214 100028
rect 101278 99958 101306 100028
rect 101266 99952 101318 99958
rect 101266 99894 101318 99900
rect 101186 99742 101260 99770
rect 100944 99680 100996 99686
rect 100772 99606 100892 99634
rect 100944 99622 100996 99628
rect 101128 99680 101180 99686
rect 101128 99622 101180 99628
rect 100760 99544 100812 99550
rect 100760 99486 100812 99492
rect 100666 98424 100722 98433
rect 100666 98359 100722 98368
rect 100574 98152 100630 98161
rect 100574 98087 100630 98096
rect 100496 95206 100616 95234
rect 100588 94602 100616 95206
rect 100404 94574 100616 94602
rect 100668 94580 100720 94586
rect 100404 94364 100432 94574
rect 100668 94522 100720 94528
rect 100404 94336 100524 94364
rect 100496 86954 100524 94336
rect 100404 86926 100524 86954
rect 100300 82340 100352 82346
rect 100300 82282 100352 82288
rect 100404 77294 100432 86926
rect 100576 82340 100628 82346
rect 100576 82282 100628 82288
rect 100404 77266 100524 77294
rect 100496 39778 100524 77266
rect 100484 39772 100536 39778
rect 100484 39714 100536 39720
rect 100588 9314 100616 82282
rect 100576 9308 100628 9314
rect 100576 9250 100628 9256
rect 100680 7818 100708 94522
rect 100772 22914 100800 99486
rect 100864 26042 100892 99606
rect 100956 94704 100984 99622
rect 101036 99408 101088 99414
rect 101036 99350 101088 99356
rect 101048 96422 101076 99350
rect 101036 96416 101088 96422
rect 101036 96358 101088 96364
rect 100956 94676 101076 94704
rect 100944 94580 100996 94586
rect 100944 94522 100996 94528
rect 100852 26036 100904 26042
rect 100852 25978 100904 25984
rect 100956 25906 100984 94522
rect 101048 94450 101076 94676
rect 101036 94444 101088 94450
rect 101036 94386 101088 94392
rect 101036 92540 101088 92546
rect 101036 92482 101088 92488
rect 100944 25900 100996 25906
rect 100944 25842 100996 25848
rect 101048 25838 101076 92482
rect 101140 25974 101168 99622
rect 101232 94858 101260 99742
rect 101370 99736 101398 100028
rect 101462 99958 101490 100028
rect 101450 99952 101502 99958
rect 101450 99894 101502 99900
rect 101554 99822 101582 100028
rect 101646 99963 101674 100028
rect 101632 99954 101688 99963
rect 101738 99958 101766 100028
rect 101830 99963 101858 100028
rect 101632 99889 101688 99898
rect 101726 99952 101778 99958
rect 101726 99894 101778 99900
rect 101816 99954 101872 99963
rect 101816 99889 101872 99898
rect 101542 99816 101594 99822
rect 101542 99758 101594 99764
rect 101922 99736 101950 100028
rect 102014 99963 102042 100028
rect 102000 99954 102056 99963
rect 102106 99958 102134 100028
rect 102198 99958 102226 100028
rect 102290 99958 102318 100028
rect 102382 99958 102410 100028
rect 102474 99958 102502 100028
rect 102566 99963 102594 100028
rect 102000 99889 102056 99898
rect 102094 99952 102146 99958
rect 102094 99894 102146 99900
rect 102186 99952 102238 99958
rect 102186 99894 102238 99900
rect 102278 99952 102330 99958
rect 102278 99894 102330 99900
rect 102370 99952 102422 99958
rect 102370 99894 102422 99900
rect 102462 99952 102514 99958
rect 102462 99894 102514 99900
rect 102552 99954 102608 99963
rect 102552 99889 102608 99898
rect 102658 99890 102686 100028
rect 102750 99963 102778 100028
rect 102736 99954 102792 99963
rect 102842 99958 102870 100028
rect 102646 99884 102698 99890
rect 102736 99889 102792 99898
rect 102830 99952 102882 99958
rect 102830 99894 102882 99900
rect 102646 99826 102698 99832
rect 102048 99816 102100 99822
rect 102048 99758 102100 99764
rect 102324 99816 102376 99822
rect 102934 99804 102962 100028
rect 103026 99822 103054 100028
rect 103118 99963 103146 100028
rect 103104 99954 103160 99963
rect 103104 99889 103160 99898
rect 102888 99793 102962 99804
rect 102324 99758 102376 99764
rect 102506 99784 102562 99793
rect 101370 99708 101444 99736
rect 101922 99708 101996 99736
rect 101416 99618 101444 99708
rect 101588 99680 101640 99686
rect 101968 99657 101996 99708
rect 101588 99622 101640 99628
rect 101678 99648 101734 99657
rect 101312 99612 101364 99618
rect 101312 99554 101364 99560
rect 101404 99612 101456 99618
rect 101404 99554 101456 99560
rect 101496 99612 101548 99618
rect 101496 99554 101548 99560
rect 101220 94852 101272 94858
rect 101220 94794 101272 94800
rect 101220 94444 101272 94450
rect 101220 94386 101272 94392
rect 101232 41138 101260 94386
rect 101324 86562 101352 99554
rect 101402 99512 101458 99521
rect 101402 99447 101458 99456
rect 101416 86630 101444 99447
rect 101508 88194 101536 99554
rect 101600 94586 101628 99622
rect 101954 99648 102010 99657
rect 101678 99583 101734 99592
rect 101864 99612 101916 99618
rect 101588 94580 101640 94586
rect 101588 94522 101640 94528
rect 101692 92546 101720 99583
rect 101954 99583 102010 99592
rect 101864 99554 101916 99560
rect 101770 98288 101826 98297
rect 101770 98223 101826 98232
rect 101784 95713 101812 98223
rect 101770 95704 101826 95713
rect 101770 95639 101826 95648
rect 101876 94790 101904 99554
rect 101956 99544 102008 99550
rect 101956 99486 102008 99492
rect 101968 97442 101996 99486
rect 102060 98394 102088 99758
rect 102336 99600 102364 99758
rect 102416 99748 102468 99754
rect 102506 99719 102562 99728
rect 102874 99784 102962 99793
rect 102930 99776 102962 99784
rect 103014 99816 103066 99822
rect 103014 99758 103066 99764
rect 102874 99719 102930 99728
rect 102416 99690 102468 99696
rect 102244 99572 102364 99600
rect 102048 98388 102100 98394
rect 102048 98330 102100 98336
rect 102046 98288 102102 98297
rect 102046 98223 102102 98232
rect 101956 97436 102008 97442
rect 101956 97378 102008 97384
rect 102060 95577 102088 98223
rect 102140 95600 102192 95606
rect 102046 95568 102102 95577
rect 102140 95542 102192 95548
rect 102046 95503 102102 95512
rect 101864 94784 101916 94790
rect 101864 94726 101916 94732
rect 101680 92540 101732 92546
rect 101680 92482 101732 92488
rect 101496 88188 101548 88194
rect 101496 88130 101548 88136
rect 101404 86624 101456 86630
rect 101404 86566 101456 86572
rect 101312 86556 101364 86562
rect 101312 86498 101364 86504
rect 101220 41132 101272 41138
rect 101220 41074 101272 41080
rect 101128 25968 101180 25974
rect 101128 25910 101180 25916
rect 101036 25832 101088 25838
rect 101036 25774 101088 25780
rect 100760 22908 100812 22914
rect 100760 22850 100812 22856
rect 102152 9178 102180 95542
rect 102244 95470 102272 99572
rect 102322 99512 102378 99521
rect 102322 99447 102378 99456
rect 102232 95464 102284 95470
rect 102232 95406 102284 95412
rect 102336 95282 102364 99447
rect 102244 95254 102364 95282
rect 102140 9172 102192 9178
rect 102140 9114 102192 9120
rect 102244 9110 102272 95254
rect 102428 91094 102456 99690
rect 102336 91066 102456 91094
rect 102336 9246 102364 91066
rect 102416 90160 102468 90166
rect 102416 90102 102468 90108
rect 102428 10742 102456 90102
rect 102520 22778 102548 99719
rect 102968 99680 103020 99686
rect 102782 99648 102838 99657
rect 102600 99612 102652 99618
rect 103210 99668 103238 100028
rect 103302 99958 103330 100028
rect 103290 99952 103342 99958
rect 103290 99894 103342 99900
rect 103394 99822 103422 100028
rect 103486 99958 103514 100028
rect 103474 99952 103526 99958
rect 103578 99929 103606 100028
rect 103474 99894 103526 99900
rect 103564 99920 103620 99929
rect 103670 99890 103698 100028
rect 103762 99958 103790 100028
rect 103854 99958 103882 100028
rect 103946 99958 103974 100028
rect 104038 99958 104066 100028
rect 104130 99958 104158 100028
rect 103750 99952 103802 99958
rect 103750 99894 103802 99900
rect 103842 99952 103894 99958
rect 103842 99894 103894 99900
rect 103934 99952 103986 99958
rect 103934 99894 103986 99900
rect 104026 99952 104078 99958
rect 104026 99894 104078 99900
rect 104118 99952 104170 99958
rect 104118 99894 104170 99900
rect 104222 99895 104250 100028
rect 103564 99855 103620 99864
rect 103658 99884 103710 99890
rect 103658 99826 103710 99832
rect 104208 99886 104264 99895
rect 103290 99816 103342 99822
rect 103288 99784 103290 99793
rect 103382 99816 103434 99822
rect 104208 99821 104264 99830
rect 103342 99784 103344 99793
rect 103382 99758 103434 99764
rect 103288 99719 103344 99728
rect 103888 99748 103940 99754
rect 104314 99736 104342 100028
rect 104406 99958 104434 100028
rect 104394 99952 104446 99958
rect 104394 99894 104446 99900
rect 104498 99890 104526 100028
rect 104590 99929 104618 100028
rect 104682 99958 104710 100028
rect 104670 99952 104722 99958
rect 104576 99920 104632 99929
rect 104486 99884 104538 99890
rect 104670 99894 104722 99900
rect 104774 99906 104802 100028
rect 104958 99963 104986 100028
rect 104944 99954 105000 99963
rect 104774 99890 104848 99906
rect 104774 99884 104860 99890
rect 104944 99889 105000 99898
rect 105050 99890 105078 100028
rect 105142 99958 105170 100028
rect 105130 99952 105182 99958
rect 105130 99894 105182 99900
rect 104774 99878 104808 99884
rect 104576 99855 104632 99864
rect 104486 99826 104538 99832
rect 104808 99826 104860 99832
rect 105038 99884 105090 99890
rect 105038 99826 105090 99832
rect 104624 99816 104676 99822
rect 104624 99758 104676 99764
rect 104990 99784 105046 99793
rect 104314 99708 104388 99736
rect 103888 99690 103940 99696
rect 103336 99680 103388 99686
rect 103210 99640 103284 99668
rect 102968 99622 103020 99628
rect 102782 99583 102838 99592
rect 102600 99554 102652 99560
rect 102612 95606 102640 99554
rect 102692 99544 102744 99550
rect 102692 99486 102744 99492
rect 102600 95600 102652 95606
rect 102600 95542 102652 95548
rect 102600 95464 102652 95470
rect 102600 95406 102652 95412
rect 102612 22846 102640 95406
rect 102704 27130 102732 99486
rect 102692 27124 102744 27130
rect 102692 27066 102744 27072
rect 102796 27062 102824 99583
rect 102876 99408 102928 99414
rect 102876 99350 102928 99356
rect 102888 27198 102916 99350
rect 102980 90166 103008 99622
rect 103256 98512 103284 99640
rect 103334 99648 103336 99657
rect 103388 99648 103390 99657
rect 103518 99648 103574 99657
rect 103334 99583 103390 99592
rect 103428 99612 103480 99618
rect 103518 99583 103574 99592
rect 103428 99554 103480 99560
rect 103336 99544 103388 99550
rect 103336 99486 103388 99492
rect 103164 98484 103284 98512
rect 103058 98288 103114 98297
rect 103058 98223 103114 98232
rect 103072 95577 103100 98223
rect 103058 95568 103114 95577
rect 103058 95503 103114 95512
rect 103164 91769 103192 98484
rect 103244 98388 103296 98394
rect 103244 98330 103296 98336
rect 103150 91760 103206 91769
rect 103150 91695 103206 91704
rect 102968 90160 103020 90166
rect 102968 90102 103020 90108
rect 103256 89282 103284 98330
rect 103348 94722 103376 99486
rect 103336 94716 103388 94722
rect 103336 94658 103388 94664
rect 103440 92818 103468 99554
rect 103532 96558 103560 99583
rect 103612 99544 103664 99550
rect 103612 99486 103664 99492
rect 103704 99544 103756 99550
rect 103704 99486 103756 99492
rect 103624 98297 103652 99486
rect 103610 98288 103666 98297
rect 103610 98223 103666 98232
rect 103612 98184 103664 98190
rect 103612 98126 103664 98132
rect 103520 96552 103572 96558
rect 103520 96494 103572 96500
rect 103520 96076 103572 96082
rect 103520 96018 103572 96024
rect 103428 92812 103480 92818
rect 103428 92754 103480 92760
rect 103244 89276 103296 89282
rect 103244 89218 103296 89224
rect 102876 27192 102928 27198
rect 102876 27134 102928 27140
rect 102784 27056 102836 27062
rect 102784 26998 102836 27004
rect 102600 22840 102652 22846
rect 102600 22782 102652 22788
rect 102508 22772 102560 22778
rect 102508 22714 102560 22720
rect 102416 10736 102468 10742
rect 102416 10678 102468 10684
rect 102324 9240 102376 9246
rect 102324 9182 102376 9188
rect 102232 9104 102284 9110
rect 102232 9046 102284 9052
rect 103532 9042 103560 96018
rect 103624 95928 103652 98126
rect 103716 96082 103744 99486
rect 103796 99476 103848 99482
rect 103796 99418 103848 99424
rect 103808 98190 103836 99418
rect 103796 98184 103848 98190
rect 103796 98126 103848 98132
rect 103900 96614 103928 99690
rect 103980 99680 104032 99686
rect 103980 99622 104032 99628
rect 104072 99680 104124 99686
rect 104072 99622 104124 99628
rect 104162 99648 104218 99657
rect 103808 96586 103928 96614
rect 103704 96076 103756 96082
rect 103704 96018 103756 96024
rect 103624 95900 103744 95928
rect 103612 95804 103664 95810
rect 103612 95746 103664 95752
rect 103624 10606 103652 95746
rect 103716 10674 103744 95900
rect 103808 26926 103836 96586
rect 103888 96552 103940 96558
rect 103888 96494 103940 96500
rect 103900 26994 103928 96494
rect 103992 28626 104020 99622
rect 104084 95656 104112 99622
rect 104162 99583 104218 99592
rect 104176 95826 104204 99583
rect 104256 99408 104308 99414
rect 104256 99350 104308 99356
rect 104268 96529 104296 99350
rect 104254 96520 104310 96529
rect 104254 96455 104310 96464
rect 104176 95798 104296 95826
rect 104360 95810 104388 99708
rect 104440 99680 104492 99686
rect 104440 99622 104492 99628
rect 104530 99648 104586 99657
rect 104268 95656 104296 95798
rect 104348 95804 104400 95810
rect 104348 95746 104400 95752
rect 104452 95713 104480 99622
rect 104530 99583 104586 99592
rect 104438 95704 104494 95713
rect 104084 95628 104204 95656
rect 104268 95628 104388 95656
rect 104438 95639 104494 95648
rect 104070 95568 104126 95577
rect 104070 95503 104126 95512
rect 104084 28694 104112 95503
rect 104072 28688 104124 28694
rect 104072 28630 104124 28636
rect 103980 28620 104032 28626
rect 103980 28562 104032 28568
rect 104176 28558 104204 95628
rect 104256 92812 104308 92818
rect 104256 92754 104308 92760
rect 104268 86494 104296 92754
rect 104256 86488 104308 86494
rect 104256 86430 104308 86436
rect 104360 86426 104388 95628
rect 104544 89214 104572 99583
rect 104636 95577 104664 99758
rect 104716 99748 104768 99754
rect 104716 99690 104768 99696
rect 104900 99748 104952 99754
rect 104990 99719 105046 99728
rect 104900 99690 104952 99696
rect 104622 95568 104678 95577
rect 104622 95503 104678 95512
rect 104728 94489 104756 99690
rect 104808 99680 104860 99686
rect 104806 99648 104808 99657
rect 104860 99648 104862 99657
rect 104806 99583 104862 99592
rect 104912 97578 104940 99690
rect 104900 97572 104952 97578
rect 104900 97514 104952 97520
rect 104900 97300 104952 97306
rect 104900 97242 104952 97248
rect 104714 94480 104770 94489
rect 104714 94415 104770 94424
rect 104532 89208 104584 89214
rect 104532 89150 104584 89156
rect 104438 87544 104494 87553
rect 104438 87479 104494 87488
rect 104348 86420 104400 86426
rect 104348 86362 104400 86368
rect 104164 28552 104216 28558
rect 104164 28494 104216 28500
rect 103888 26988 103940 26994
rect 103888 26930 103940 26936
rect 103796 26920 103848 26926
rect 103796 26862 103848 26868
rect 103704 10668 103756 10674
rect 103704 10610 103756 10616
rect 103612 10600 103664 10606
rect 103612 10542 103664 10548
rect 103520 9036 103572 9042
rect 103520 8978 103572 8984
rect 100668 7812 100720 7818
rect 100668 7754 100720 7760
rect 100392 5500 100444 5506
rect 100392 5442 100444 5448
rect 100116 5296 100168 5302
rect 100116 5238 100168 5244
rect 100024 3392 100076 3398
rect 100024 3334 100076 3340
rect 100404 480 100432 5442
rect 103704 5228 103756 5234
rect 103704 5170 103756 5176
rect 102600 3732 102652 3738
rect 102600 3674 102652 3680
rect 101496 3392 101548 3398
rect 101496 3334 101548 3340
rect 101508 480 101536 3334
rect 102612 480 102640 3674
rect 103716 480 103744 5170
rect 104452 3738 104480 87479
rect 104912 5234 104940 97242
rect 105004 95742 105032 99719
rect 105084 99612 105136 99618
rect 105084 99554 105136 99560
rect 105096 96014 105124 99554
rect 105234 99532 105262 100028
rect 105326 99958 105354 100028
rect 105314 99952 105366 99958
rect 105314 99894 105366 99900
rect 105418 99890 105446 100028
rect 105510 99958 105538 100028
rect 105498 99952 105550 99958
rect 105602 99929 105630 100028
rect 105498 99894 105550 99900
rect 105588 99920 105644 99929
rect 105406 99884 105458 99890
rect 105588 99855 105644 99864
rect 105406 99826 105458 99832
rect 105694 99736 105722 100028
rect 105648 99708 105722 99736
rect 105544 99680 105596 99686
rect 105544 99622 105596 99628
rect 105452 99544 105504 99550
rect 105188 99504 105262 99532
rect 105372 99504 105452 99532
rect 105188 97034 105216 99504
rect 105266 98288 105322 98297
rect 105266 98223 105322 98232
rect 105176 97028 105228 97034
rect 105176 96970 105228 96976
rect 105176 96892 105228 96898
rect 105176 96834 105228 96840
rect 105084 96008 105136 96014
rect 105084 95950 105136 95956
rect 105084 95872 105136 95878
rect 105084 95814 105136 95820
rect 104992 95736 105044 95742
rect 104992 95678 105044 95684
rect 104992 95600 105044 95606
rect 104992 95542 105044 95548
rect 105004 10470 105032 95542
rect 105096 10538 105124 95814
rect 105188 95606 105216 96834
rect 105176 95600 105228 95606
rect 105176 95542 105228 95548
rect 105176 93968 105228 93974
rect 105176 93910 105228 93916
rect 105084 10532 105136 10538
rect 105084 10474 105136 10480
rect 104992 10464 105044 10470
rect 104992 10406 105044 10412
rect 105188 10402 105216 93910
rect 105280 28354 105308 98223
rect 105372 95878 105400 99504
rect 105452 99486 105504 99492
rect 105556 97306 105584 99622
rect 105544 97300 105596 97306
rect 105544 97242 105596 97248
rect 105452 97028 105504 97034
rect 105452 96970 105504 96976
rect 105360 95872 105412 95878
rect 105360 95814 105412 95820
rect 105360 95736 105412 95742
rect 105360 95678 105412 95684
rect 105372 28490 105400 95678
rect 105360 28484 105412 28490
rect 105360 28426 105412 28432
rect 105464 28422 105492 96970
rect 105648 96898 105676 99708
rect 105786 99668 105814 100028
rect 105740 99640 105814 99668
rect 105636 96892 105688 96898
rect 105636 96834 105688 96840
rect 105740 96778 105768 99640
rect 105878 99600 105906 100028
rect 105970 99890 105998 100028
rect 106062 99963 106090 100028
rect 106048 99954 106104 99963
rect 105958 99884 106010 99890
rect 106048 99889 106104 99898
rect 106154 99890 106182 100028
rect 106246 99958 106274 100028
rect 106338 99958 106366 100028
rect 106234 99952 106286 99958
rect 106234 99894 106286 99900
rect 106326 99952 106378 99958
rect 106326 99894 106378 99900
rect 105958 99826 106010 99832
rect 106142 99884 106194 99890
rect 106142 99826 106194 99832
rect 106430 99822 106458 100028
rect 106522 99958 106550 100028
rect 106510 99952 106562 99958
rect 106510 99894 106562 99900
rect 106418 99816 106470 99822
rect 106418 99758 106470 99764
rect 106004 99748 106056 99754
rect 106004 99690 106056 99696
rect 106280 99748 106332 99754
rect 106614 99736 106642 100028
rect 106706 99958 106734 100028
rect 106694 99952 106746 99958
rect 106694 99894 106746 99900
rect 106280 99690 106332 99696
rect 106568 99708 106642 99736
rect 106798 99736 106826 100028
rect 106890 99958 106918 100028
rect 106982 99958 107010 100028
rect 107074 99958 107102 100028
rect 106878 99952 106930 99958
rect 106878 99894 106930 99900
rect 106970 99952 107022 99958
rect 106970 99894 107022 99900
rect 107062 99952 107114 99958
rect 107062 99894 107114 99900
rect 106924 99816 106976 99822
rect 106924 99758 106976 99764
rect 106798 99708 106872 99736
rect 105556 96750 105768 96778
rect 105832 99572 105906 99600
rect 105556 41002 105584 96750
rect 105832 96614 105860 99572
rect 106016 99498 106044 99690
rect 106096 99680 106148 99686
rect 106096 99622 106148 99628
rect 106188 99680 106240 99686
rect 106188 99622 106240 99628
rect 105648 96586 105860 96614
rect 105924 99470 106044 99498
rect 105648 41070 105676 96586
rect 105728 96008 105780 96014
rect 105728 95950 105780 95956
rect 105740 89146 105768 95950
rect 105924 93974 105952 99470
rect 106004 99408 106056 99414
rect 106004 99350 106056 99356
rect 106016 94654 106044 99350
rect 106108 96257 106136 99622
rect 106200 97510 106228 99622
rect 106188 97504 106240 97510
rect 106188 97446 106240 97452
rect 106292 96626 106320 99690
rect 106372 99612 106424 99618
rect 106372 99554 106424 99560
rect 106280 96620 106332 96626
rect 106280 96562 106332 96568
rect 106094 96248 106150 96257
rect 106384 96234 106412 99554
rect 106464 99476 106516 99482
rect 106464 99418 106516 99424
rect 106476 96762 106504 99418
rect 106464 96756 106516 96762
rect 106464 96698 106516 96704
rect 106462 96656 106518 96665
rect 106462 96591 106518 96600
rect 106094 96183 106150 96192
rect 106292 96206 106412 96234
rect 106292 96014 106320 96206
rect 106372 96076 106424 96082
rect 106372 96018 106424 96024
rect 106280 96008 106332 96014
rect 106280 95950 106332 95956
rect 106280 95872 106332 95878
rect 106280 95814 106332 95820
rect 106004 94648 106056 94654
rect 106004 94590 106056 94596
rect 105912 93968 105964 93974
rect 105912 93910 105964 93916
rect 105728 89140 105780 89146
rect 105728 89082 105780 89088
rect 105636 41064 105688 41070
rect 105636 41006 105688 41012
rect 105544 40996 105596 41002
rect 105544 40938 105596 40944
rect 105452 28416 105504 28422
rect 105452 28358 105504 28364
rect 105268 28348 105320 28354
rect 105268 28290 105320 28296
rect 106292 12102 106320 95814
rect 106384 12170 106412 96018
rect 106476 29850 106504 96591
rect 106568 29986 106596 99708
rect 106648 99612 106700 99618
rect 106648 99554 106700 99560
rect 106556 29980 106608 29986
rect 106556 29922 106608 29928
rect 106660 29918 106688 99554
rect 106740 99544 106792 99550
rect 106740 99486 106792 99492
rect 106752 96801 106780 99486
rect 106738 96792 106794 96801
rect 106738 96727 106794 96736
rect 106740 96620 106792 96626
rect 106740 96562 106792 96568
rect 106752 30122 106780 96562
rect 106844 96150 106872 99708
rect 106832 96144 106884 96150
rect 106832 96086 106884 96092
rect 106832 96008 106884 96014
rect 106832 95950 106884 95956
rect 106740 30116 106792 30122
rect 106740 30058 106792 30064
rect 106844 30054 106872 95950
rect 106936 31414 106964 99758
rect 107016 99748 107068 99754
rect 107166 99736 107194 100028
rect 107016 99690 107068 99696
rect 107120 99708 107194 99736
rect 107028 96082 107056 99690
rect 107120 99374 107148 99708
rect 107258 99668 107286 100028
rect 107442 99940 107470 100028
rect 107396 99929 107470 99940
rect 107534 99929 107562 100028
rect 107626 99958 107654 100028
rect 107718 99958 107746 100028
rect 107614 99952 107666 99958
rect 107382 99920 107470 99929
rect 107438 99912 107470 99920
rect 107520 99920 107576 99929
rect 107382 99855 107438 99864
rect 107614 99894 107666 99900
rect 107706 99952 107758 99958
rect 107706 99894 107758 99900
rect 107520 99855 107576 99864
rect 107660 99816 107712 99822
rect 107566 99784 107622 99793
rect 107476 99748 107528 99754
rect 107810 99804 107838 100028
rect 107902 99963 107930 100028
rect 107888 99954 107944 99963
rect 107994 99958 108022 100028
rect 107888 99889 107944 99898
rect 107982 99952 108034 99958
rect 107982 99894 108034 99900
rect 107810 99776 107884 99804
rect 107660 99758 107712 99764
rect 107566 99719 107622 99728
rect 107476 99690 107528 99696
rect 107258 99640 107332 99668
rect 107488 99657 107516 99690
rect 107120 99346 107240 99374
rect 107108 96756 107160 96762
rect 107108 96698 107160 96704
rect 107016 96076 107068 96082
rect 107016 96018 107068 96024
rect 107016 95940 107068 95946
rect 107016 95882 107068 95888
rect 107028 82278 107056 95882
rect 107120 90438 107148 96698
rect 107212 95878 107240 99346
rect 107304 96393 107332 99640
rect 107474 99648 107530 99657
rect 107384 99612 107436 99618
rect 107474 99583 107530 99592
rect 107384 99554 107436 99560
rect 107290 96384 107346 96393
rect 107290 96319 107346 96328
rect 107396 96150 107424 99554
rect 107474 99512 107530 99521
rect 107474 99447 107530 99456
rect 107384 96144 107436 96150
rect 107384 96086 107436 96092
rect 107200 95872 107252 95878
rect 107200 95814 107252 95820
rect 107488 94926 107516 99447
rect 107580 96257 107608 99719
rect 107672 99668 107700 99758
rect 107856 99736 107884 99776
rect 108086 99736 108114 100028
rect 107856 99708 107930 99736
rect 107672 99640 107792 99668
rect 107658 99512 107714 99521
rect 107658 99447 107714 99456
rect 107566 96248 107622 96257
rect 107566 96183 107622 96192
rect 107476 94920 107528 94926
rect 107476 94862 107528 94868
rect 107108 90432 107160 90438
rect 107108 90374 107160 90380
rect 107016 82272 107068 82278
rect 107016 82214 107068 82220
rect 106924 31408 106976 31414
rect 106924 31350 106976 31356
rect 106832 30048 106884 30054
rect 106832 29990 106884 29996
rect 106648 29912 106700 29918
rect 106648 29854 106700 29860
rect 106464 29844 106516 29850
rect 106464 29786 106516 29792
rect 106372 12164 106424 12170
rect 106372 12106 106424 12112
rect 106280 12096 106332 12102
rect 106280 12038 106332 12044
rect 107672 12034 107700 99447
rect 107764 95606 107792 99640
rect 107902 99634 107930 99708
rect 107856 99606 107930 99634
rect 108040 99708 108114 99736
rect 108178 99736 108206 100028
rect 108270 99963 108298 100028
rect 108256 99954 108312 99963
rect 108362 99958 108390 100028
rect 108256 99889 108312 99898
rect 108350 99952 108402 99958
rect 108350 99894 108402 99900
rect 108454 99804 108482 100028
rect 108546 99958 108574 100028
rect 108638 99963 108666 100028
rect 108534 99952 108586 99958
rect 108534 99894 108586 99900
rect 108624 99954 108680 99963
rect 108624 99889 108680 99898
rect 108408 99793 108482 99804
rect 108394 99784 108482 99793
rect 108178 99708 108252 99736
rect 108450 99776 108482 99784
rect 108394 99719 108450 99728
rect 107752 95600 107804 95606
rect 107752 95542 107804 95548
rect 107750 95432 107806 95441
rect 107750 95367 107806 95376
rect 107660 12028 107712 12034
rect 107660 11970 107712 11976
rect 107764 11898 107792 95367
rect 107856 94178 107884 99606
rect 107936 96144 107988 96150
rect 107936 96086 107988 96092
rect 107844 94172 107896 94178
rect 107844 94114 107896 94120
rect 107844 94036 107896 94042
rect 107844 93978 107896 93984
rect 107856 11966 107884 93978
rect 107948 90386 107976 96086
rect 108040 93498 108068 99708
rect 108120 99612 108172 99618
rect 108120 99554 108172 99560
rect 108028 93492 108080 93498
rect 108028 93434 108080 93440
rect 108132 91094 108160 99554
rect 108224 94042 108252 99708
rect 108730 99668 108758 100028
rect 108822 99895 108850 100028
rect 108808 99886 108864 99895
rect 108808 99821 108864 99830
rect 108810 99748 108862 99754
rect 108914 99736 108942 100028
rect 109006 99822 109034 100028
rect 109098 99958 109126 100028
rect 109086 99952 109138 99958
rect 109086 99894 109138 99900
rect 108994 99816 109046 99822
rect 109190 99770 109218 100028
rect 108994 99758 109046 99764
rect 108862 99708 108942 99736
rect 109144 99742 109218 99770
rect 109282 99770 109310 100028
rect 109374 99890 109402 100028
rect 109466 99929 109494 100028
rect 109452 99920 109508 99929
rect 109362 99884 109414 99890
rect 109452 99855 109508 99864
rect 109362 99826 109414 99832
rect 109558 99804 109586 100028
rect 109512 99776 109586 99804
rect 109282 99742 109356 99770
rect 108810 99690 108862 99696
rect 108684 99657 108758 99668
rect 108302 99648 108358 99657
rect 108302 99583 108358 99592
rect 108670 99648 108758 99657
rect 108726 99640 108758 99648
rect 109040 99680 109092 99686
rect 109040 99622 109092 99628
rect 108670 99583 108726 99592
rect 108948 99612 109000 99618
rect 108212 94036 108264 94042
rect 108212 93978 108264 93984
rect 108132 91066 108252 91094
rect 107948 90358 108160 90386
rect 107936 90296 107988 90302
rect 107936 90238 107988 90244
rect 107948 13462 107976 90238
rect 108028 90228 108080 90234
rect 108028 90170 108080 90176
rect 107936 13456 107988 13462
rect 107936 13398 107988 13404
rect 108040 13394 108068 90170
rect 108132 29782 108160 90358
rect 108120 29776 108172 29782
rect 108120 29718 108172 29724
rect 108224 29714 108252 91066
rect 108316 90302 108344 99583
rect 108948 99554 109000 99560
rect 108396 99544 108448 99550
rect 108396 99486 108448 99492
rect 108672 99544 108724 99550
rect 108672 99486 108724 99492
rect 108762 99512 108818 99521
rect 108304 90296 108356 90302
rect 108304 90238 108356 90244
rect 108304 90160 108356 90166
rect 108304 90102 108356 90108
rect 108316 31346 108344 90102
rect 108408 32842 108436 99486
rect 108488 99476 108540 99482
rect 108488 99418 108540 99424
rect 108500 99374 108528 99418
rect 108500 99346 108620 99374
rect 108488 94172 108540 94178
rect 108488 94114 108540 94120
rect 108500 90166 108528 94114
rect 108592 90234 108620 99346
rect 108684 96257 108712 99486
rect 108762 99447 108818 99456
rect 108776 96665 108804 99447
rect 108960 99374 108988 99554
rect 108868 99346 108988 99374
rect 108762 96656 108818 96665
rect 108762 96591 108818 96600
rect 108670 96248 108726 96257
rect 108670 96183 108726 96192
rect 108764 95600 108816 95606
rect 108764 95542 108816 95548
rect 108580 90228 108632 90234
rect 108580 90170 108632 90176
rect 108488 90160 108540 90166
rect 108488 90102 108540 90108
rect 108776 85134 108804 95542
rect 108868 94450 108896 99346
rect 109052 96150 109080 99622
rect 109144 96626 109172 99742
rect 109132 96620 109184 96626
rect 109132 96562 109184 96568
rect 109328 96234 109356 99742
rect 109512 96234 109540 99776
rect 109650 99736 109678 100028
rect 109144 96206 109356 96234
rect 109420 96206 109540 96234
rect 109604 99708 109678 99736
rect 109742 99736 109770 100028
rect 109834 99958 109862 100028
rect 109926 100026 109954 100028
rect 109914 100020 109966 100026
rect 109914 99962 109966 99968
rect 110018 99958 110046 100028
rect 110110 99958 110138 100028
rect 109822 99952 109874 99958
rect 109822 99894 109874 99900
rect 110006 99952 110058 99958
rect 110006 99894 110058 99900
rect 110098 99952 110150 99958
rect 110202 99929 110230 100028
rect 110098 99894 110150 99900
rect 110188 99920 110244 99929
rect 110294 99890 110322 100028
rect 110386 99890 110414 100028
rect 110478 99958 110506 100028
rect 110466 99952 110518 99958
rect 110466 99894 110518 99900
rect 110188 99855 110244 99864
rect 110282 99884 110334 99890
rect 110282 99826 110334 99832
rect 110374 99884 110426 99890
rect 110374 99826 110426 99832
rect 110570 99822 110598 100028
rect 110558 99816 110610 99822
rect 110662 99793 110690 100028
rect 110754 99804 110782 100028
rect 110846 99958 110874 100028
rect 110834 99952 110886 99958
rect 110834 99894 110886 99900
rect 110558 99758 110610 99764
rect 110648 99784 110704 99793
rect 110052 99748 110104 99754
rect 109742 99708 109816 99736
rect 109040 96144 109092 96150
rect 109040 96086 109092 96092
rect 108948 94512 109000 94518
rect 108948 94454 109000 94460
rect 108856 94444 108908 94450
rect 108856 94386 108908 94392
rect 108960 92474 108988 94454
rect 108960 92446 109080 92474
rect 108764 85128 108816 85134
rect 108764 85070 108816 85076
rect 108396 32836 108448 32842
rect 108396 32778 108448 32784
rect 108304 31340 108356 31346
rect 108304 31282 108356 31288
rect 108212 29708 108264 29714
rect 108212 29650 108264 29656
rect 108028 13388 108080 13394
rect 108028 13330 108080 13336
rect 107844 11960 107896 11966
rect 107844 11902 107896 11908
rect 107752 11892 107804 11898
rect 107752 11834 107804 11840
rect 109052 11830 109080 92446
rect 109144 13326 109172 96206
rect 109224 96076 109276 96082
rect 109224 96018 109276 96024
rect 109132 13320 109184 13326
rect 109132 13262 109184 13268
rect 109236 13190 109264 96018
rect 109420 95962 109448 96206
rect 109500 96144 109552 96150
rect 109500 96086 109552 96092
rect 109328 95934 109448 95962
rect 109328 13258 109356 95934
rect 109408 95668 109460 95674
rect 109408 95610 109460 95616
rect 109420 14822 109448 95610
rect 109512 31278 109540 96086
rect 109604 94586 109632 99708
rect 109684 99476 109736 99482
rect 109684 99418 109736 99424
rect 109592 94580 109644 94586
rect 109592 94522 109644 94528
rect 109592 94444 109644 94450
rect 109592 94386 109644 94392
rect 109604 39710 109632 94386
rect 109696 83502 109724 99418
rect 109788 93362 109816 99708
rect 110052 99690 110104 99696
rect 110144 99748 110196 99754
rect 110144 99690 110196 99696
rect 110420 99748 110472 99754
rect 110754 99776 110828 99804
rect 110648 99719 110704 99728
rect 110420 99690 110472 99696
rect 109868 99680 109920 99686
rect 109868 99622 109920 99628
rect 109880 96082 109908 99622
rect 109960 99544 110012 99550
rect 109960 99486 110012 99492
rect 109868 96076 109920 96082
rect 109868 96018 109920 96024
rect 109972 95674 110000 99486
rect 110064 96257 110092 99690
rect 110050 96248 110106 96257
rect 110050 96183 110106 96192
rect 109960 95668 110012 95674
rect 109960 95610 110012 95616
rect 110156 93401 110184 99690
rect 110236 99680 110288 99686
rect 110236 99622 110288 99628
rect 110248 96801 110276 99622
rect 110326 98152 110382 98161
rect 110326 98087 110382 98096
rect 110234 96792 110290 96801
rect 110234 96727 110290 96736
rect 110236 96620 110288 96626
rect 110236 96562 110288 96568
rect 110248 95130 110276 96562
rect 110236 95124 110288 95130
rect 110236 95066 110288 95072
rect 110340 93770 110368 98087
rect 110432 97306 110460 99690
rect 110512 99680 110564 99686
rect 110512 99622 110564 99628
rect 110602 99648 110658 99657
rect 110420 97300 110472 97306
rect 110420 97242 110472 97248
rect 110524 97050 110552 99622
rect 110602 99583 110658 99592
rect 110616 97170 110644 99583
rect 110696 99544 110748 99550
rect 110696 99486 110748 99492
rect 110604 97164 110656 97170
rect 110604 97106 110656 97112
rect 110524 97022 110644 97050
rect 110418 96520 110474 96529
rect 110418 96455 110474 96464
rect 110328 93764 110380 93770
rect 110328 93706 110380 93712
rect 110142 93392 110198 93401
rect 109776 93356 109828 93362
rect 110142 93327 110198 93336
rect 109776 93298 109828 93304
rect 109684 83496 109736 83502
rect 109684 83438 109736 83444
rect 109592 39704 109644 39710
rect 109592 39646 109644 39652
rect 109500 31272 109552 31278
rect 109500 31214 109552 31220
rect 109408 14816 109460 14822
rect 109408 14758 109460 14764
rect 109316 13252 109368 13258
rect 109316 13194 109368 13200
rect 109224 13184 109276 13190
rect 109224 13126 109276 13132
rect 110432 13122 110460 96455
rect 110512 95600 110564 95606
rect 110512 95542 110564 95548
rect 110524 14754 110552 95542
rect 110616 24206 110644 97022
rect 110708 28286 110736 99486
rect 110800 31142 110828 99776
rect 110938 99736 110966 100028
rect 111030 99958 111058 100028
rect 111122 99958 111150 100028
rect 111018 99952 111070 99958
rect 111018 99894 111070 99900
rect 111110 99952 111162 99958
rect 111214 99929 111242 100028
rect 111110 99894 111162 99900
rect 111200 99920 111256 99929
rect 111200 99855 111256 99864
rect 111156 99816 111208 99822
rect 111156 99758 111208 99764
rect 111306 99770 111334 100028
rect 111398 99963 111426 100028
rect 111384 99954 111440 99963
rect 111384 99889 111440 99898
rect 111490 99890 111518 100028
rect 111582 99958 111610 100028
rect 111570 99952 111622 99958
rect 111570 99894 111622 99900
rect 111674 99890 111702 100028
rect 111766 99929 111794 100028
rect 111752 99920 111808 99929
rect 111478 99884 111530 99890
rect 111478 99826 111530 99832
rect 111662 99884 111714 99890
rect 111858 99890 111886 100028
rect 111752 99855 111808 99864
rect 111846 99884 111898 99890
rect 111662 99826 111714 99832
rect 111846 99826 111898 99832
rect 111706 99784 111762 99793
rect 110938 99708 111012 99736
rect 110880 99544 110932 99550
rect 110880 99486 110932 99492
rect 110788 31136 110840 31142
rect 110788 31078 110840 31084
rect 110892 31074 110920 99486
rect 110984 98122 111012 99708
rect 111064 99612 111116 99618
rect 111064 99554 111116 99560
rect 110972 98116 111024 98122
rect 110972 98058 111024 98064
rect 110972 97980 111024 97986
rect 110972 97922 111024 97928
rect 110984 34270 111012 97922
rect 111076 34338 111104 99554
rect 111168 97986 111196 99758
rect 111306 99742 111380 99770
rect 111352 99618 111380 99742
rect 111432 99748 111484 99754
rect 111950 99770 111978 100028
rect 112042 99958 112070 100028
rect 112030 99952 112082 99958
rect 112030 99894 112082 99900
rect 112134 99770 112162 100028
rect 111762 99742 111840 99770
rect 111706 99719 111762 99728
rect 111432 99690 111484 99696
rect 111340 99612 111392 99618
rect 111340 99554 111392 99560
rect 111338 99512 111394 99521
rect 111338 99447 111394 99456
rect 111156 97980 111208 97986
rect 111156 97922 111208 97928
rect 111156 97164 111208 97170
rect 111156 97106 111208 97112
rect 111168 88126 111196 97106
rect 111352 93430 111380 99447
rect 111444 95577 111472 99690
rect 111616 99680 111668 99686
rect 111616 99622 111668 99628
rect 111524 99612 111576 99618
rect 111524 99554 111576 99560
rect 111536 95606 111564 99554
rect 111628 99385 111656 99622
rect 111708 99612 111760 99618
rect 111708 99554 111760 99560
rect 111614 99376 111670 99385
rect 111614 99311 111670 99320
rect 111616 99272 111668 99278
rect 111616 99214 111668 99220
rect 111628 96830 111656 99214
rect 111616 96824 111668 96830
rect 111616 96766 111668 96772
rect 111720 96393 111748 99554
rect 111706 96384 111762 96393
rect 111706 96319 111762 96328
rect 111524 95600 111576 95606
rect 111430 95568 111486 95577
rect 111524 95542 111576 95548
rect 111430 95503 111486 95512
rect 111812 94738 111840 99742
rect 111720 94710 111840 94738
rect 111904 99742 111978 99770
rect 112088 99742 112162 99770
rect 111720 94178 111748 94710
rect 111800 94580 111852 94586
rect 111800 94522 111852 94528
rect 111708 94172 111760 94178
rect 111708 94114 111760 94120
rect 111524 93764 111576 93770
rect 111524 93706 111576 93712
rect 111340 93424 111392 93430
rect 111340 93366 111392 93372
rect 111156 88120 111208 88126
rect 111156 88062 111208 88068
rect 111536 84194 111564 93706
rect 111444 84166 111564 84194
rect 111064 34332 111116 34338
rect 111064 34274 111116 34280
rect 110972 34264 111024 34270
rect 110972 34206 111024 34212
rect 111444 31210 111472 84166
rect 111432 31204 111484 31210
rect 111432 31146 111484 31152
rect 110880 31068 110932 31074
rect 110880 31010 110932 31016
rect 110696 28280 110748 28286
rect 110696 28222 110748 28228
rect 110604 24200 110656 24206
rect 110604 24142 110656 24148
rect 110604 21412 110656 21418
rect 110604 21354 110656 21360
rect 110616 16574 110644 21354
rect 110616 16546 111472 16574
rect 110512 14748 110564 14754
rect 110512 14690 110564 14696
rect 110420 13116 110472 13122
rect 110420 13058 110472 13064
rect 109040 11824 109092 11830
rect 109040 11766 109092 11772
rect 105176 10396 105228 10402
rect 105176 10338 105228 10344
rect 106188 6384 106240 6390
rect 106188 6326 106240 6332
rect 104900 5228 104952 5234
rect 104900 5170 104952 5176
rect 106200 4010 106228 6326
rect 107016 5092 107068 5098
rect 107016 5034 107068 5040
rect 106188 4004 106240 4010
rect 106188 3946 106240 3952
rect 104808 3936 104860 3942
rect 104808 3878 104860 3884
rect 104440 3732 104492 3738
rect 104440 3674 104492 3680
rect 104820 480 104848 3878
rect 105910 3496 105966 3505
rect 105910 3431 105966 3440
rect 105924 480 105952 3431
rect 107028 480 107056 5034
rect 108120 5024 108172 5030
rect 108120 4966 108172 4972
rect 108132 480 108160 4966
rect 110328 4956 110380 4962
rect 110328 4898 110380 4904
rect 109224 3800 109276 3806
rect 109224 3742 109276 3748
rect 109236 480 109264 3742
rect 110340 480 110368 4898
rect 111444 480 111472 16546
rect 111812 14686 111840 94522
rect 111904 25770 111932 99742
rect 111984 99680 112036 99686
rect 112088 99657 112116 99742
rect 112226 99668 112254 100028
rect 112318 99890 112346 100028
rect 112306 99884 112358 99890
rect 112306 99826 112358 99832
rect 112410 99770 112438 100028
rect 111984 99622 112036 99628
rect 112074 99648 112130 99657
rect 111996 99498 112024 99622
rect 112074 99583 112130 99592
rect 112180 99640 112254 99668
rect 112364 99742 112438 99770
rect 111996 99470 112116 99498
rect 111984 99408 112036 99414
rect 111984 99350 112036 99356
rect 111996 94586 112024 99350
rect 112088 94586 112116 99470
rect 111984 94580 112036 94586
rect 111984 94522 112036 94528
rect 112076 94580 112128 94586
rect 112076 94522 112128 94528
rect 112180 94466 112208 99640
rect 112258 99376 112314 99385
rect 112258 99311 112314 99320
rect 111996 94438 112208 94466
rect 111892 25764 111944 25770
rect 111892 25706 111944 25712
rect 111996 25702 112024 94438
rect 112168 94376 112220 94382
rect 112168 94318 112220 94324
rect 112076 94308 112128 94314
rect 112076 94250 112128 94256
rect 111984 25696 112036 25702
rect 111984 25638 112036 25644
rect 112088 25634 112116 94250
rect 112180 32638 112208 94318
rect 112272 32774 112300 99311
rect 112260 32768 112312 32774
rect 112260 32710 112312 32716
rect 112364 32706 112392 99742
rect 112502 99668 112530 100028
rect 112686 99906 112714 100028
rect 112456 99640 112530 99668
rect 112640 99878 112714 99906
rect 112456 94314 112484 99640
rect 112640 99498 112668 99878
rect 112778 99804 112806 100028
rect 112548 99470 112668 99498
rect 112732 99776 112806 99804
rect 112548 94382 112576 99470
rect 112628 99408 112680 99414
rect 112628 99350 112680 99356
rect 112536 94376 112588 94382
rect 112536 94318 112588 94324
rect 112444 94308 112496 94314
rect 112444 94250 112496 94256
rect 112536 94240 112588 94246
rect 112536 94182 112588 94188
rect 112444 94172 112496 94178
rect 112444 94114 112496 94120
rect 112456 39642 112484 94114
rect 112548 85066 112576 94182
rect 112536 85060 112588 85066
rect 112536 85002 112588 85008
rect 112640 84998 112668 99350
rect 112732 96801 112760 99776
rect 112870 99668 112898 100028
rect 112824 99640 112898 99668
rect 112962 99668 112990 100028
rect 113054 99770 113082 100028
rect 113146 99890 113174 100028
rect 113134 99884 113186 99890
rect 113134 99826 113186 99832
rect 113238 99770 113266 100028
rect 113330 99929 113358 100028
rect 113316 99920 113372 99929
rect 113316 99855 113372 99864
rect 113422 99770 113450 100028
rect 113514 99890 113542 100028
rect 113502 99884 113554 99890
rect 113502 99826 113554 99832
rect 113606 99770 113634 100028
rect 113698 99958 113726 100028
rect 113686 99952 113738 99958
rect 113686 99894 113738 99900
rect 113790 99770 113818 100028
rect 113882 100026 113910 100028
rect 113870 100020 113922 100026
rect 113870 99962 113922 99968
rect 113974 99906 114002 100028
rect 113054 99742 113128 99770
rect 112962 99640 113036 99668
rect 112824 96937 112852 99640
rect 113008 99498 113036 99640
rect 112916 99470 113036 99498
rect 112810 96928 112866 96937
rect 112810 96863 112866 96872
rect 112812 96824 112864 96830
rect 112718 96792 112774 96801
rect 112812 96766 112864 96772
rect 112718 96727 112774 96736
rect 112824 93294 112852 96766
rect 112916 96665 112944 99470
rect 113100 99374 113128 99742
rect 113008 99346 113128 99374
rect 113192 99742 113266 99770
rect 113376 99742 113450 99770
rect 113560 99742 113634 99770
rect 113744 99742 113818 99770
rect 113928 99878 114002 99906
rect 113008 97073 113036 99346
rect 113088 97980 113140 97986
rect 113088 97922 113140 97928
rect 112994 97064 113050 97073
rect 112994 96999 113050 97008
rect 113100 96830 113128 97922
rect 113088 96824 113140 96830
rect 113088 96766 113140 96772
rect 112902 96656 112958 96665
rect 112902 96591 112958 96600
rect 113192 94738 113220 99742
rect 113272 99680 113324 99686
rect 113272 99622 113324 99628
rect 113100 94710 113220 94738
rect 113100 94382 113128 94710
rect 113284 94602 113312 99622
rect 113192 94574 113312 94602
rect 113088 94376 113140 94382
rect 113088 94318 113140 94324
rect 112812 93288 112864 93294
rect 112812 93230 112864 93236
rect 112628 84992 112680 84998
rect 112628 84934 112680 84940
rect 112444 39636 112496 39642
rect 112444 39578 112496 39584
rect 112352 32700 112404 32706
rect 112352 32642 112404 32648
rect 112168 32632 112220 32638
rect 112168 32574 112220 32580
rect 112076 25628 112128 25634
rect 112076 25570 112128 25576
rect 111800 14680 111852 14686
rect 111800 14622 111852 14628
rect 113192 14550 113220 94574
rect 113272 94444 113324 94450
rect 113272 94386 113324 94392
rect 113180 14544 113232 14550
rect 113180 14486 113232 14492
rect 113284 14482 113312 94386
rect 113376 14618 113404 99742
rect 113456 99612 113508 99618
rect 113456 99554 113508 99560
rect 113468 95062 113496 99554
rect 113456 95056 113508 95062
rect 113456 94998 113508 95004
rect 113560 94602 113588 99742
rect 113640 99680 113692 99686
rect 113640 99622 113692 99628
rect 113468 94574 113588 94602
rect 113468 25566 113496 94574
rect 113548 94512 113600 94518
rect 113548 94454 113600 94460
rect 113560 32434 113588 94454
rect 113652 32502 113680 99622
rect 113744 94518 113772 99742
rect 113928 99686 113956 99878
rect 114066 99770 114094 100028
rect 114158 99958 114186 100028
rect 114146 99952 114198 99958
rect 114146 99894 114198 99900
rect 114250 99770 114278 100028
rect 114342 99793 114370 100028
rect 114020 99742 114094 99770
rect 114204 99742 114278 99770
rect 114328 99784 114384 99793
rect 113824 99680 113876 99686
rect 113824 99622 113876 99628
rect 113916 99680 113968 99686
rect 113916 99622 113968 99628
rect 113836 97986 113864 99622
rect 113914 99512 113970 99521
rect 113914 99447 113970 99456
rect 113824 97980 113876 97986
rect 113824 97922 113876 97928
rect 113928 97617 113956 99447
rect 113914 97608 113970 97617
rect 113824 97572 113876 97578
rect 113914 97543 113970 97552
rect 113824 97514 113876 97520
rect 113836 96762 113864 97514
rect 113916 97504 113968 97510
rect 113916 97446 113968 97452
rect 113824 96756 113876 96762
rect 113824 96698 113876 96704
rect 113824 95056 113876 95062
rect 113824 94998 113876 95004
rect 113732 94512 113784 94518
rect 113732 94454 113784 94460
rect 113732 94376 113784 94382
rect 113732 94318 113784 94324
rect 113744 32570 113772 94318
rect 113836 82210 113864 94998
rect 113928 90506 113956 97446
rect 114020 96665 114048 99742
rect 114100 99680 114152 99686
rect 114100 99622 114152 99628
rect 114006 96656 114062 96665
rect 114006 96591 114062 96600
rect 114112 94450 114140 99622
rect 114204 96801 114232 99742
rect 114328 99719 114384 99728
rect 114434 99736 114462 100028
rect 114526 99929 114554 100028
rect 114512 99920 114568 99929
rect 114512 99855 114568 99864
rect 114618 99770 114646 100028
rect 114710 99958 114738 100028
rect 114698 99952 114750 99958
rect 114698 99894 114750 99900
rect 114572 99742 114646 99770
rect 114434 99708 114508 99736
rect 114480 99600 114508 99708
rect 114388 99572 114508 99600
rect 114284 98116 114336 98122
rect 114284 98058 114336 98064
rect 114190 96792 114246 96801
rect 114190 96727 114246 96736
rect 114100 94444 114152 94450
rect 114100 94386 114152 94392
rect 114296 92002 114324 98058
rect 114388 96937 114416 99572
rect 114468 99476 114520 99482
rect 114468 99418 114520 99424
rect 114374 96928 114430 96937
rect 114374 96863 114430 96872
rect 114374 96792 114430 96801
rect 114374 96727 114430 96736
rect 114388 93226 114416 96727
rect 114480 94314 114508 99418
rect 114572 94450 114600 99742
rect 114802 99736 114830 100028
rect 114894 99958 114922 100028
rect 114882 99952 114934 99958
rect 114882 99894 114934 99900
rect 114986 99890 115014 100028
rect 114974 99884 115026 99890
rect 114974 99826 115026 99832
rect 115078 99770 115106 100028
rect 115170 99958 115198 100028
rect 115158 99952 115210 99958
rect 115158 99894 115210 99900
rect 115262 99770 115290 100028
rect 115354 99958 115382 100028
rect 115446 99958 115474 100028
rect 115342 99952 115394 99958
rect 115342 99894 115394 99900
rect 115434 99952 115486 99958
rect 115434 99894 115486 99900
rect 115538 99770 115566 100028
rect 115032 99759 115106 99770
rect 114756 99708 114830 99736
rect 115018 99750 115106 99759
rect 114650 99648 114706 99657
rect 114650 99583 114706 99592
rect 114560 94444 114612 94450
rect 114560 94386 114612 94392
rect 114468 94308 114520 94314
rect 114468 94250 114520 94256
rect 114376 93220 114428 93226
rect 114376 93162 114428 93168
rect 114284 91996 114336 92002
rect 114284 91938 114336 91944
rect 113916 90500 113968 90506
rect 113916 90442 113968 90448
rect 114560 90024 114612 90030
rect 114560 89966 114612 89972
rect 113824 82204 113876 82210
rect 113824 82146 113876 82152
rect 113732 32564 113784 32570
rect 113732 32506 113784 32512
rect 113640 32496 113692 32502
rect 113640 32438 113692 32444
rect 113548 32428 113600 32434
rect 113548 32370 113600 32376
rect 113456 25560 113508 25566
rect 113456 25502 113508 25508
rect 114572 16114 114600 89966
rect 114664 16250 114692 99583
rect 114756 99532 114784 99708
rect 115074 99742 115106 99750
rect 115216 99742 115290 99770
rect 115354 99742 115566 99770
rect 115018 99685 115074 99694
rect 115112 99680 115164 99686
rect 115112 99622 115164 99628
rect 115020 99612 115072 99618
rect 115020 99554 115072 99560
rect 114928 99544 114980 99550
rect 114756 99504 114876 99532
rect 114744 99340 114796 99346
rect 114744 99282 114796 99288
rect 114756 95044 114784 99282
rect 114848 95198 114876 99504
rect 114928 99486 114980 99492
rect 114940 96966 114968 99486
rect 114928 96960 114980 96966
rect 114928 96902 114980 96908
rect 114928 96824 114980 96830
rect 114928 96766 114980 96772
rect 114940 96150 114968 96766
rect 114928 96144 114980 96150
rect 114928 96086 114980 96092
rect 114928 96008 114980 96014
rect 114928 95950 114980 95956
rect 114836 95192 114888 95198
rect 114836 95134 114888 95140
rect 114756 95016 114876 95044
rect 114744 94376 114796 94382
rect 114744 94318 114796 94324
rect 114652 16244 114704 16250
rect 114652 16186 114704 16192
rect 114756 16182 114784 94318
rect 114848 19038 114876 95016
rect 114940 34066 114968 95950
rect 115032 34134 115060 99554
rect 115124 96014 115152 99622
rect 115216 99550 115244 99742
rect 115354 99668 115382 99742
rect 115308 99640 115382 99668
rect 115480 99680 115532 99686
rect 115204 99544 115256 99550
rect 115204 99486 115256 99492
rect 115202 99388 115258 99397
rect 115202 99323 115258 99332
rect 115112 96008 115164 96014
rect 115112 95950 115164 95956
rect 115216 94602 115244 99323
rect 115308 94738 115336 99640
rect 115630 99668 115658 100028
rect 115722 99822 115750 100028
rect 115710 99816 115762 99822
rect 115710 99758 115762 99764
rect 115480 99622 115532 99628
rect 115584 99640 115658 99668
rect 115388 99544 115440 99550
rect 115388 99486 115440 99492
rect 115400 95282 115428 99486
rect 115492 95418 115520 99622
rect 115584 96665 115612 99640
rect 115814 99634 115842 100028
rect 115906 99958 115934 100028
rect 115998 99958 116026 100028
rect 116090 99958 116118 100028
rect 116182 99963 116210 100028
rect 115894 99952 115946 99958
rect 115894 99894 115946 99900
rect 115986 99952 116038 99958
rect 115986 99894 116038 99900
rect 116078 99952 116130 99958
rect 116078 99894 116130 99900
rect 116168 99954 116224 99963
rect 116168 99889 116224 99898
rect 116274 99890 116302 100028
rect 116366 99963 116394 100028
rect 116352 99954 116408 99963
rect 116458 99958 116486 100028
rect 116262 99884 116314 99890
rect 116352 99889 116408 99898
rect 116446 99952 116498 99958
rect 116550 99929 116578 100028
rect 116642 99958 116670 100028
rect 116734 99958 116762 100028
rect 116826 99958 116854 100028
rect 116630 99952 116682 99958
rect 116446 99894 116498 99900
rect 116536 99920 116592 99929
rect 116630 99894 116682 99900
rect 116722 99952 116774 99958
rect 116722 99894 116774 99900
rect 116814 99952 116866 99958
rect 116814 99894 116866 99900
rect 116536 99855 116592 99864
rect 116262 99826 116314 99832
rect 116492 99816 116544 99822
rect 116398 99784 116454 99793
rect 116124 99748 116176 99754
rect 116492 99758 116544 99764
rect 116918 99770 116946 100028
rect 117010 99958 117038 100028
rect 117102 99963 117130 100028
rect 116998 99952 117050 99958
rect 116998 99894 117050 99900
rect 117088 99954 117144 99963
rect 117088 99889 117144 99898
rect 117194 99770 117222 100028
rect 117286 99890 117314 100028
rect 117378 99958 117406 100028
rect 117470 99958 117498 100028
rect 117562 99958 117590 100028
rect 117366 99952 117418 99958
rect 117366 99894 117418 99900
rect 117458 99952 117510 99958
rect 117458 99894 117510 99900
rect 117550 99952 117602 99958
rect 117746 99906 117774 100028
rect 117838 99958 117866 100028
rect 117930 99958 117958 100028
rect 117550 99894 117602 99900
rect 117274 99884 117326 99890
rect 117274 99826 117326 99832
rect 117700 99878 117774 99906
rect 117826 99952 117878 99958
rect 117826 99894 117878 99900
rect 117918 99952 117970 99958
rect 117918 99894 117970 99900
rect 118022 99890 118050 100028
rect 118010 99884 118062 99890
rect 116398 99719 116454 99728
rect 116124 99690 116176 99696
rect 115768 99606 115842 99634
rect 116032 99612 116084 99618
rect 115664 99544 115716 99550
rect 115664 99486 115716 99492
rect 115676 96801 115704 99486
rect 115768 96830 115796 99606
rect 116136 99600 116164 99690
rect 116308 99680 116360 99686
rect 116308 99622 116360 99628
rect 116136 99572 116256 99600
rect 116032 99554 116084 99560
rect 115848 99544 115900 99550
rect 115848 99486 115900 99492
rect 115940 99544 115992 99550
rect 115940 99486 115992 99492
rect 115756 96824 115808 96830
rect 115662 96792 115718 96801
rect 115756 96766 115808 96772
rect 115662 96727 115718 96736
rect 115570 96656 115626 96665
rect 115570 96591 115626 96600
rect 115756 96144 115808 96150
rect 115756 96086 115808 96092
rect 115492 95390 115704 95418
rect 115400 95254 115612 95282
rect 115480 95192 115532 95198
rect 115480 95134 115532 95140
rect 115308 94710 115428 94738
rect 115216 94574 115336 94602
rect 115204 94512 115256 94518
rect 115204 94454 115256 94460
rect 115112 94444 115164 94450
rect 115112 94386 115164 94392
rect 115124 34202 115152 94386
rect 115216 35494 115244 94454
rect 115308 87990 115336 94574
rect 115400 94518 115428 94710
rect 115388 94512 115440 94518
rect 115388 94454 115440 94460
rect 115492 89714 115520 95134
rect 115584 94382 115612 95254
rect 115572 94376 115624 94382
rect 115572 94318 115624 94324
rect 115676 90030 115704 95390
rect 115768 93158 115796 96086
rect 115860 95402 115888 99486
rect 115848 95396 115900 95402
rect 115848 95338 115900 95344
rect 115848 95124 115900 95130
rect 115848 95066 115900 95072
rect 115860 94518 115888 95066
rect 115848 94512 115900 94518
rect 115848 94454 115900 94460
rect 115756 93152 115808 93158
rect 115756 93094 115808 93100
rect 115664 90024 115716 90030
rect 115664 89966 115716 89972
rect 115400 89686 115520 89714
rect 115400 89078 115428 89686
rect 115388 89072 115440 89078
rect 115388 89014 115440 89020
rect 115296 87984 115348 87990
rect 115296 87926 115348 87932
rect 115388 87644 115440 87650
rect 115388 87586 115440 87592
rect 115204 35488 115256 35494
rect 115204 35430 115256 35436
rect 115112 34196 115164 34202
rect 115112 34138 115164 34144
rect 115020 34128 115072 34134
rect 115020 34070 115072 34076
rect 114928 34060 114980 34066
rect 114928 34002 114980 34008
rect 114836 19032 114888 19038
rect 114836 18974 114888 18980
rect 114744 16176 114796 16182
rect 114744 16118 114796 16124
rect 114560 16108 114612 16114
rect 114560 16050 114612 16056
rect 113364 14612 113416 14618
rect 113364 14554 113416 14560
rect 113272 14476 113324 14482
rect 113272 14418 113324 14424
rect 114744 6316 114796 6322
rect 114744 6258 114796 6264
rect 113640 6248 113692 6254
rect 113640 6190 113692 6196
rect 112536 3596 112588 3602
rect 112536 3538 112588 3544
rect 112548 480 112576 3538
rect 113652 480 113680 6190
rect 114756 480 114784 6258
rect 115400 3942 115428 87586
rect 115952 16046 115980 99486
rect 116044 95062 116072 99554
rect 116122 99512 116178 99521
rect 116122 99447 116178 99456
rect 116032 95056 116084 95062
rect 116032 94998 116084 95004
rect 116032 94580 116084 94586
rect 116032 94522 116084 94528
rect 116044 33998 116072 94522
rect 116032 33992 116084 33998
rect 116032 33934 116084 33940
rect 116136 33930 116164 99447
rect 116228 38010 116256 99572
rect 116320 94586 116348 99622
rect 116412 97594 116440 99719
rect 116504 99346 116532 99758
rect 116584 99748 116636 99754
rect 116918 99742 116992 99770
rect 117194 99742 117268 99770
rect 117700 99754 117728 99878
rect 118010 99826 118062 99832
rect 116584 99690 116636 99696
rect 116492 99340 116544 99346
rect 116492 99282 116544 99288
rect 116412 97566 116532 97594
rect 116400 97368 116452 97374
rect 116400 97310 116452 97316
rect 116412 96558 116440 97310
rect 116400 96552 116452 96558
rect 116400 96494 116452 96500
rect 116400 95056 116452 95062
rect 116400 94998 116452 95004
rect 116308 94580 116360 94586
rect 116308 94522 116360 94528
rect 116308 94444 116360 94450
rect 116308 94386 116360 94392
rect 116216 38004 116268 38010
rect 116216 37946 116268 37952
rect 116320 37942 116348 94386
rect 116412 40934 116440 94998
rect 116504 84930 116532 97566
rect 116596 86358 116624 99690
rect 116860 99680 116912 99686
rect 116860 99622 116912 99628
rect 116768 99612 116820 99618
rect 116768 99554 116820 99560
rect 116676 99136 116728 99142
rect 116676 99078 116728 99084
rect 116688 89010 116716 99078
rect 116780 97481 116808 99554
rect 116766 97472 116822 97481
rect 116766 97407 116822 97416
rect 116872 96614 116900 99622
rect 116780 96586 116900 96614
rect 116780 94450 116808 96586
rect 116860 96552 116912 96558
rect 116860 96494 116912 96500
rect 116768 94444 116820 94450
rect 116768 94386 116820 94392
rect 116872 92274 116900 96494
rect 116964 95810 116992 99742
rect 117136 99680 117188 99686
rect 117240 99657 117268 99742
rect 117504 99748 117556 99754
rect 117504 99690 117556 99696
rect 117688 99748 117740 99754
rect 118114 99736 118142 100028
rect 118206 99890 118234 100028
rect 118298 99929 118326 100028
rect 118390 99958 118418 100028
rect 118482 99963 118510 100028
rect 118378 99952 118430 99958
rect 118284 99920 118340 99929
rect 118194 99884 118246 99890
rect 118378 99894 118430 99900
rect 118468 99954 118524 99963
rect 118468 99889 118524 99898
rect 118284 99855 118340 99864
rect 118194 99826 118246 99832
rect 118238 99784 118294 99793
rect 118114 99708 118188 99736
rect 118238 99719 118240 99728
rect 117688 99690 117740 99696
rect 117136 99622 117188 99628
rect 117226 99648 117282 99657
rect 117148 98326 117176 99622
rect 117516 99634 117544 99690
rect 117872 99680 117924 99686
rect 117226 99583 117282 99592
rect 117412 99612 117464 99618
rect 117516 99606 117636 99634
rect 117872 99622 117924 99628
rect 117412 99554 117464 99560
rect 117226 99512 117282 99521
rect 117226 99447 117228 99456
rect 117280 99447 117282 99456
rect 117320 99476 117372 99482
rect 117228 99418 117280 99424
rect 117320 99418 117372 99424
rect 117136 98320 117188 98326
rect 117136 98262 117188 98268
rect 117044 96824 117096 96830
rect 117044 96766 117096 96772
rect 116952 95804 117004 95810
rect 116952 95746 117004 95752
rect 116860 92268 116912 92274
rect 116860 92210 116912 92216
rect 117056 89714 117084 96766
rect 117332 94466 117360 99418
rect 117424 94602 117452 99554
rect 117504 99544 117556 99550
rect 117504 99486 117556 99492
rect 117516 96150 117544 99486
rect 117608 98410 117636 99606
rect 117780 99544 117832 99550
rect 117780 99486 117832 99492
rect 117608 98382 117728 98410
rect 117596 98320 117648 98326
rect 117596 98262 117648 98268
rect 117504 96144 117556 96150
rect 117504 96086 117556 96092
rect 117608 94976 117636 98262
rect 117700 96558 117728 98382
rect 117688 96552 117740 96558
rect 117688 96494 117740 96500
rect 117688 96144 117740 96150
rect 117688 96086 117740 96092
rect 117516 94948 117636 94976
rect 117516 94738 117544 94948
rect 117516 94710 117636 94738
rect 117424 94574 117544 94602
rect 117332 94438 117452 94466
rect 117320 94376 117372 94382
rect 117320 94318 117372 94324
rect 116964 89686 117084 89714
rect 116676 89004 116728 89010
rect 116676 88946 116728 88952
rect 116584 86352 116636 86358
rect 116584 86294 116636 86300
rect 116492 84924 116544 84930
rect 116492 84866 116544 84872
rect 116400 40928 116452 40934
rect 116400 40870 116452 40876
rect 116964 38078 116992 89686
rect 116952 38072 117004 38078
rect 116952 38014 117004 38020
rect 116308 37936 116360 37942
rect 116308 37878 116360 37884
rect 116124 33924 116176 33930
rect 116124 33866 116176 33872
rect 117332 33862 117360 94318
rect 117424 35358 117452 94438
rect 117516 35426 117544 94574
rect 117608 39574 117636 94710
rect 117700 84862 117728 96086
rect 117792 86290 117820 99486
rect 117884 94382 117912 99622
rect 117964 99612 118016 99618
rect 118160 99600 118188 99708
rect 118292 99719 118294 99728
rect 118574 99736 118602 100028
rect 118666 99958 118694 100028
rect 118654 99952 118706 99958
rect 118654 99894 118706 99900
rect 118758 99890 118786 100028
rect 118746 99884 118798 99890
rect 118746 99826 118798 99832
rect 118850 99770 118878 100028
rect 118942 99963 118970 100028
rect 118928 99954 118984 99963
rect 118928 99889 118984 99898
rect 118850 99742 118924 99770
rect 118574 99708 118648 99736
rect 118240 99690 118292 99696
rect 118424 99612 118476 99618
rect 118160 99572 118280 99600
rect 117964 99554 118016 99560
rect 117976 97986 118004 99554
rect 117964 97980 118016 97986
rect 117964 97922 118016 97928
rect 118148 97572 118200 97578
rect 118148 97514 118200 97520
rect 118160 97102 118188 97514
rect 118148 97096 118200 97102
rect 118252 97073 118280 99572
rect 118424 99554 118476 99560
rect 118332 99476 118384 99482
rect 118332 99418 118384 99424
rect 118148 97038 118200 97044
rect 118238 97064 118294 97073
rect 118344 97050 118372 99418
rect 118436 97209 118464 99554
rect 118620 97238 118648 99708
rect 118698 99648 118754 99657
rect 118698 99583 118754 99592
rect 118608 97232 118660 97238
rect 118422 97200 118478 97209
rect 118608 97174 118660 97180
rect 118422 97135 118478 97144
rect 118344 97022 118648 97050
rect 118238 96999 118294 97008
rect 118330 96928 118386 96937
rect 118330 96863 118386 96872
rect 118344 96506 118372 96863
rect 118516 96824 118568 96830
rect 118516 96766 118568 96772
rect 118344 96478 118464 96506
rect 118148 95396 118200 95402
rect 118148 95338 118200 95344
rect 117872 94376 117924 94382
rect 117872 94318 117924 94324
rect 118160 89714 118188 95338
rect 118332 94444 118384 94450
rect 118332 94386 118384 94392
rect 118160 89686 118280 89714
rect 117780 86284 117832 86290
rect 117780 86226 117832 86232
rect 117688 84856 117740 84862
rect 117688 84798 117740 84804
rect 117596 39568 117648 39574
rect 117596 39510 117648 39516
rect 118252 36582 118280 89686
rect 118344 38146 118372 94386
rect 118436 87922 118464 96478
rect 118528 94450 118556 96766
rect 118516 94444 118568 94450
rect 118516 94386 118568 94392
rect 118620 91934 118648 97022
rect 118608 91928 118660 91934
rect 118608 91870 118660 91876
rect 118424 87916 118476 87922
rect 118424 87858 118476 87864
rect 118332 38140 118384 38146
rect 118332 38082 118384 38088
rect 118240 36576 118292 36582
rect 118240 36518 118292 36524
rect 117504 35420 117556 35426
rect 117504 35362 117556 35368
rect 117412 35352 117464 35358
rect 117412 35294 117464 35300
rect 117320 33856 117372 33862
rect 117320 33798 117372 33804
rect 118712 17542 118740 99583
rect 118792 99544 118844 99550
rect 118792 99486 118844 99492
rect 118804 96966 118832 99486
rect 118792 96960 118844 96966
rect 118792 96902 118844 96908
rect 118896 96898 118924 99742
rect 119034 99736 119062 100028
rect 119126 99804 119154 100028
rect 119218 99958 119246 100028
rect 119206 99952 119258 99958
rect 119206 99894 119258 99900
rect 119310 99822 119338 100028
rect 119298 99816 119350 99822
rect 119126 99776 119200 99804
rect 119034 99708 119108 99736
rect 118976 99612 119028 99618
rect 118976 99554 119028 99560
rect 118988 97442 119016 99554
rect 118976 97436 119028 97442
rect 118976 97378 119028 97384
rect 118976 97300 119028 97306
rect 118976 97242 119028 97248
rect 118884 96892 118936 96898
rect 118884 96834 118936 96840
rect 118792 96824 118844 96830
rect 118792 96766 118844 96772
rect 118700 17536 118752 17542
rect 118700 17478 118752 17484
rect 118804 17474 118832 96766
rect 118884 96620 118936 96626
rect 118884 96562 118936 96568
rect 118896 18834 118924 96562
rect 118988 24138 119016 97242
rect 119080 40798 119108 99708
rect 119172 97170 119200 99776
rect 119298 99758 119350 99764
rect 119402 99634 119430 100028
rect 119494 99958 119522 100028
rect 119586 99958 119614 100028
rect 119678 99958 119706 100028
rect 119482 99952 119534 99958
rect 119482 99894 119534 99900
rect 119574 99952 119626 99958
rect 119574 99894 119626 99900
rect 119666 99952 119718 99958
rect 119770 99929 119798 100028
rect 119666 99894 119718 99900
rect 119756 99920 119812 99929
rect 119862 99890 119890 100028
rect 119954 99890 119982 100028
rect 120046 99958 120074 100028
rect 120138 99958 120166 100028
rect 120034 99952 120086 99958
rect 120034 99894 120086 99900
rect 120126 99952 120178 99958
rect 120126 99894 120178 99900
rect 119756 99855 119812 99864
rect 119850 99884 119902 99890
rect 119850 99826 119902 99832
rect 119942 99884 119994 99890
rect 119942 99826 119994 99832
rect 119528 99816 119580 99822
rect 119620 99816 119672 99822
rect 119528 99758 119580 99764
rect 119618 99784 119620 99793
rect 119712 99816 119764 99822
rect 119672 99784 119674 99793
rect 119356 99606 119430 99634
rect 119356 99498 119384 99606
rect 119264 99470 119384 99498
rect 119436 99476 119488 99482
rect 119160 97164 119212 97170
rect 119160 97106 119212 97112
rect 119160 96960 119212 96966
rect 119160 96902 119212 96908
rect 119172 40866 119200 96902
rect 119160 40860 119212 40866
rect 119160 40802 119212 40808
rect 119068 40792 119120 40798
rect 119068 40734 119120 40740
rect 119264 40730 119292 99470
rect 119436 99418 119488 99424
rect 119344 97436 119396 97442
rect 119344 97378 119396 97384
rect 119356 91866 119384 97378
rect 119448 96830 119476 99418
rect 119540 97016 119568 99758
rect 119712 99758 119764 99764
rect 120078 99784 120134 99793
rect 119618 99719 119674 99728
rect 119620 99680 119672 99686
rect 119620 99622 119672 99628
rect 119632 97306 119660 99622
rect 119724 97306 119752 99758
rect 119804 99748 119856 99754
rect 120078 99719 120134 99728
rect 120230 99736 120258 100028
rect 120322 99804 120350 100028
rect 120414 99963 120442 100028
rect 120400 99954 120456 99963
rect 120506 99958 120534 100028
rect 120598 99958 120626 100028
rect 120690 99958 120718 100028
rect 120782 99963 120810 100028
rect 120400 99889 120456 99898
rect 120494 99952 120546 99958
rect 120494 99894 120546 99900
rect 120586 99952 120638 99958
rect 120586 99894 120638 99900
rect 120678 99952 120730 99958
rect 120678 99894 120730 99900
rect 120768 99954 120824 99963
rect 120768 99889 120824 99898
rect 120724 99816 120776 99822
rect 120322 99776 120396 99804
rect 120368 99736 120396 99776
rect 120724 99758 120776 99764
rect 120874 99770 120902 100028
rect 120966 99958 120994 100028
rect 121058 99963 121086 100028
rect 120954 99952 121006 99958
rect 120954 99894 121006 99900
rect 121044 99954 121100 99963
rect 121044 99889 121100 99898
rect 121150 99804 121178 100028
rect 121242 99822 121270 100028
rect 121426 99958 121454 100028
rect 121518 99963 121546 100028
rect 121414 99952 121466 99958
rect 121414 99894 121466 99900
rect 121504 99954 121560 99963
rect 121504 99889 121560 99898
rect 121702 99895 121730 100028
rect 121688 99886 121744 99895
rect 121104 99776 121178 99804
rect 121230 99816 121282 99822
rect 121688 99821 121744 99830
rect 121104 99770 121132 99776
rect 120540 99748 120592 99754
rect 119804 99690 119856 99696
rect 119620 97300 119672 97306
rect 119620 97242 119672 97248
rect 119712 97300 119764 97306
rect 119712 97242 119764 97248
rect 119816 97209 119844 99690
rect 119896 99680 119948 99686
rect 119896 99622 119948 99628
rect 119802 97200 119858 97209
rect 119802 97135 119858 97144
rect 119804 97096 119856 97102
rect 119804 97038 119856 97044
rect 119540 96988 119660 97016
rect 119528 96892 119580 96898
rect 119528 96834 119580 96840
rect 119436 96824 119488 96830
rect 119436 96766 119488 96772
rect 119540 93838 119568 96834
rect 119632 96626 119660 96988
rect 119712 96756 119764 96762
rect 119712 96698 119764 96704
rect 119620 96620 119672 96626
rect 119620 96562 119672 96568
rect 119528 93832 119580 93838
rect 119528 93774 119580 93780
rect 119344 91860 119396 91866
rect 119344 91802 119396 91808
rect 119724 90574 119752 96698
rect 119712 90568 119764 90574
rect 119712 90510 119764 90516
rect 119344 90364 119396 90370
rect 119344 90306 119396 90312
rect 119252 40724 119304 40730
rect 119252 40666 119304 40672
rect 118976 24132 119028 24138
rect 118976 24074 119028 24080
rect 118884 18828 118936 18834
rect 118884 18770 118936 18776
rect 118792 17468 118844 17474
rect 118792 17410 118844 17416
rect 115940 16040 115992 16046
rect 115940 15982 115992 15988
rect 116952 6180 117004 6186
rect 116952 6122 117004 6128
rect 115388 3936 115440 3942
rect 115388 3878 115440 3884
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 115860 480 115888 3470
rect 116964 480 116992 6122
rect 119160 4888 119212 4894
rect 119160 4830 119212 4836
rect 118056 3460 118108 3466
rect 118056 3402 118108 3408
rect 118068 480 118096 3402
rect 119172 480 119200 4830
rect 119356 3806 119384 90306
rect 119816 89350 119844 97038
rect 119908 96121 119936 99622
rect 120092 98598 120120 99719
rect 120230 99708 120304 99736
rect 120368 99708 120442 99736
rect 120172 99612 120224 99618
rect 120172 99554 120224 99560
rect 120080 98592 120132 98598
rect 120080 98534 120132 98540
rect 120080 97368 120132 97374
rect 120080 97310 120132 97316
rect 119894 96112 119950 96121
rect 119894 96047 119950 96056
rect 120092 89714 120120 97310
rect 120184 94178 120212 99554
rect 120172 94172 120224 94178
rect 120172 94114 120224 94120
rect 120276 93854 120304 99708
rect 120414 99634 120442 99708
rect 120540 99690 120592 99696
rect 120632 99748 120684 99754
rect 120632 99690 120684 99696
rect 120368 99606 120442 99634
rect 120368 96762 120396 99606
rect 120446 99512 120502 99521
rect 120446 99447 120502 99456
rect 120356 96756 120408 96762
rect 120356 96698 120408 96704
rect 120276 93826 120396 93854
rect 120264 91792 120316 91798
rect 120264 91734 120316 91740
rect 120092 89686 120212 89714
rect 119804 89344 119856 89350
rect 119804 89286 119856 89292
rect 120184 5166 120212 89686
rect 120276 16574 120304 91734
rect 120368 17406 120396 93826
rect 120460 18766 120488 99447
rect 120552 29646 120580 99690
rect 120644 97050 120672 99690
rect 120736 97374 120764 99758
rect 120874 99742 120948 99770
rect 120816 99680 120868 99686
rect 120816 99622 120868 99628
rect 120724 97368 120776 97374
rect 120724 97310 120776 97316
rect 120828 97050 120856 99622
rect 120920 97152 120948 99742
rect 121058 99742 121132 99770
rect 121230 99758 121282 99764
rect 121058 99634 121086 99742
rect 121794 99736 121822 100028
rect 121886 99890 121914 100028
rect 121874 99884 121926 99890
rect 121874 99826 121926 99832
rect 121978 99770 122006 100028
rect 122070 99929 122098 100028
rect 122056 99920 122112 99929
rect 122056 99855 122112 99864
rect 121932 99742 122006 99770
rect 121794 99708 121868 99736
rect 121184 99680 121236 99686
rect 121058 99606 121132 99634
rect 121184 99622 121236 99628
rect 121552 99680 121604 99686
rect 121552 99622 121604 99628
rect 121642 99648 121698 99657
rect 121000 99476 121052 99482
rect 121000 99418 121052 99424
rect 121012 97345 121040 99418
rect 120998 97336 121054 97345
rect 120998 97271 121054 97280
rect 121104 97209 121132 99606
rect 121090 97200 121146 97209
rect 120920 97124 121040 97152
rect 121090 97135 121146 97144
rect 120644 97022 120764 97050
rect 120828 97022 120948 97050
rect 120630 96928 120686 96937
rect 120630 96863 120686 96872
rect 120644 33794 120672 96863
rect 120736 35290 120764 97022
rect 120816 96960 120868 96966
rect 120816 96902 120868 96908
rect 120828 39506 120856 96902
rect 120920 90370 120948 97022
rect 121012 96966 121040 97124
rect 121092 97028 121144 97034
rect 121092 96970 121144 96976
rect 121000 96960 121052 96966
rect 121000 96902 121052 96908
rect 121104 92070 121132 96970
rect 121196 96937 121224 99622
rect 121460 99612 121512 99618
rect 121460 99554 121512 99560
rect 121368 98592 121420 98598
rect 121368 98534 121420 98540
rect 121380 97578 121408 98534
rect 121368 97572 121420 97578
rect 121368 97514 121420 97520
rect 121182 96928 121238 96937
rect 121182 96863 121238 96872
rect 121368 96688 121420 96694
rect 121368 96630 121420 96636
rect 121276 94172 121328 94178
rect 121276 94114 121328 94120
rect 121092 92064 121144 92070
rect 121092 92006 121144 92012
rect 120908 90364 120960 90370
rect 120908 90306 120960 90312
rect 120816 39500 120868 39506
rect 120816 39442 120868 39448
rect 120724 35284 120776 35290
rect 120724 35226 120776 35232
rect 120632 33788 120684 33794
rect 120632 33730 120684 33736
rect 120540 29640 120592 29646
rect 120540 29582 120592 29588
rect 120448 18760 120500 18766
rect 120448 18702 120500 18708
rect 120356 17400 120408 17406
rect 120356 17342 120408 17348
rect 120276 16546 121224 16574
rect 120172 5160 120224 5166
rect 120172 5102 120224 5108
rect 120264 4820 120316 4826
rect 120264 4762 120316 4768
rect 119344 3800 119396 3806
rect 119344 3742 119396 3748
rect 120276 480 120304 4762
rect 121196 3482 121224 16546
rect 121288 3602 121316 94114
rect 121380 92342 121408 96630
rect 121472 95198 121500 99554
rect 121564 95985 121592 99622
rect 121642 99583 121698 99592
rect 121550 95976 121606 95985
rect 121550 95911 121606 95920
rect 121552 95396 121604 95402
rect 121552 95338 121604 95344
rect 121460 95192 121512 95198
rect 121460 95134 121512 95140
rect 121368 92336 121420 92342
rect 121368 92278 121420 92284
rect 121276 3596 121328 3602
rect 121276 3538 121328 3544
rect 121196 3454 121408 3482
rect 121564 3466 121592 95338
rect 121656 94994 121684 99583
rect 121736 99544 121788 99550
rect 121736 99486 121788 99492
rect 121644 94988 121696 94994
rect 121644 94930 121696 94936
rect 121644 94308 121696 94314
rect 121644 94250 121696 94256
rect 121656 5098 121684 94250
rect 121748 17270 121776 99486
rect 121840 95282 121868 99708
rect 121932 95402 121960 99742
rect 122162 99736 122190 100028
rect 122254 99958 122282 100028
rect 122346 99958 122374 100028
rect 122242 99952 122294 99958
rect 122242 99894 122294 99900
rect 122334 99952 122386 99958
rect 122334 99894 122386 99900
rect 122438 99793 122466 100028
rect 122530 99929 122558 100028
rect 122516 99920 122572 99929
rect 122516 99855 122572 99864
rect 122116 99708 122190 99736
rect 122424 99784 122480 99793
rect 122622 99770 122650 100028
rect 122714 99958 122742 100028
rect 122806 100026 122834 100028
rect 122794 100020 122846 100026
rect 122794 99962 122846 99968
rect 122702 99952 122754 99958
rect 122702 99894 122754 99900
rect 122898 99770 122926 100028
rect 122424 99719 122480 99728
rect 122576 99742 122650 99770
rect 122852 99742 122926 99770
rect 122990 99770 123018 100028
rect 123082 99890 123110 100028
rect 123070 99884 123122 99890
rect 123070 99826 123122 99832
rect 123174 99770 123202 100028
rect 123266 99958 123294 100028
rect 123254 99952 123306 99958
rect 123254 99894 123306 99900
rect 123358 99804 123386 100028
rect 123450 99958 123478 100028
rect 123542 99958 123570 100028
rect 123438 99952 123490 99958
rect 123438 99894 123490 99900
rect 123530 99952 123582 99958
rect 123530 99894 123582 99900
rect 123358 99776 123524 99804
rect 122990 99742 123064 99770
rect 123174 99742 123248 99770
rect 122116 99600 122144 99708
rect 122380 99680 122432 99686
rect 122024 99572 122144 99600
rect 122194 99648 122250 99657
rect 122380 99622 122432 99628
rect 122194 99583 122250 99592
rect 122288 99612 122340 99618
rect 122024 96150 122052 99572
rect 122102 99512 122158 99521
rect 122102 99447 122158 99456
rect 122012 96144 122064 96150
rect 122012 96086 122064 96092
rect 121920 95396 121972 95402
rect 121920 95338 121972 95344
rect 121840 95254 122052 95282
rect 121828 95192 121880 95198
rect 121828 95134 121880 95140
rect 121840 17338 121868 95134
rect 121920 94444 121972 94450
rect 121920 94386 121972 94392
rect 121932 20194 121960 94386
rect 122024 20330 122052 95254
rect 122116 20398 122144 99447
rect 122104 20392 122156 20398
rect 122104 20334 122156 20340
rect 122012 20324 122064 20330
rect 122012 20266 122064 20272
rect 122208 20262 122236 99583
rect 122288 99554 122340 99560
rect 122300 94450 122328 99554
rect 122288 94444 122340 94450
rect 122288 94386 122340 94392
rect 122392 94314 122420 99622
rect 122576 98433 122604 99742
rect 122656 99544 122708 99550
rect 122656 99486 122708 99492
rect 122562 98424 122618 98433
rect 122562 98359 122618 98368
rect 122668 96801 122696 99486
rect 122748 99476 122800 99482
rect 122748 99418 122800 99424
rect 122760 97442 122788 99418
rect 122748 97436 122800 97442
rect 122748 97378 122800 97384
rect 122654 96792 122710 96801
rect 122654 96727 122710 96736
rect 122472 95804 122524 95810
rect 122472 95746 122524 95752
rect 122380 94308 122432 94314
rect 122380 94250 122432 94256
rect 122484 80782 122512 95746
rect 122564 94988 122616 94994
rect 122564 94930 122616 94936
rect 122472 80776 122524 80782
rect 122472 80718 122524 80724
rect 122196 20256 122248 20262
rect 122196 20198 122248 20204
rect 121920 20188 121972 20194
rect 121920 20130 121972 20136
rect 121828 17332 121880 17338
rect 121828 17274 121880 17280
rect 121736 17264 121788 17270
rect 121736 17206 121788 17212
rect 121644 5092 121696 5098
rect 121644 5034 121696 5040
rect 122470 4856 122526 4865
rect 122470 4791 122526 4800
rect 121380 480 121408 3454
rect 121552 3460 121604 3466
rect 121552 3402 121604 3408
rect 122484 480 122512 4791
rect 122576 3534 122604 94930
rect 122852 94738 122880 99742
rect 122932 99680 122984 99686
rect 122932 99622 122984 99628
rect 122760 94710 122880 94738
rect 122760 94314 122788 94710
rect 122944 94602 122972 99622
rect 122852 94574 122972 94602
rect 122748 94308 122800 94314
rect 122748 94250 122800 94256
rect 122852 5030 122880 94574
rect 122932 94444 122984 94450
rect 122932 94386 122984 94392
rect 122944 6390 122972 94386
rect 123036 94382 123064 99742
rect 123116 99612 123168 99618
rect 123116 99554 123168 99560
rect 123024 94376 123076 94382
rect 123024 94318 123076 94324
rect 123024 94240 123076 94246
rect 123024 94182 123076 94188
rect 123036 18698 123064 94182
rect 123128 21554 123156 99554
rect 123220 21622 123248 99742
rect 123300 99680 123352 99686
rect 123300 99622 123352 99628
rect 123312 94994 123340 99622
rect 123392 99476 123444 99482
rect 123392 99418 123444 99424
rect 123300 94988 123352 94994
rect 123300 94930 123352 94936
rect 123404 94466 123432 99418
rect 123496 95146 123524 99776
rect 123634 99770 123662 100028
rect 123726 99890 123754 100028
rect 123714 99884 123766 99890
rect 123714 99826 123766 99832
rect 123818 99770 123846 100028
rect 123910 99929 123938 100028
rect 124002 99958 124030 100028
rect 124094 99958 124122 100028
rect 123990 99952 124042 99958
rect 123896 99920 123952 99929
rect 123990 99894 124042 99900
rect 124082 99952 124134 99958
rect 124082 99894 124134 99900
rect 124186 99890 124214 100028
rect 124278 99929 124306 100028
rect 124264 99920 124320 99929
rect 123896 99855 123952 99864
rect 124174 99884 124226 99890
rect 124370 99890 124398 100028
rect 124264 99855 124320 99864
rect 124358 99884 124410 99890
rect 124174 99826 124226 99832
rect 124358 99826 124410 99832
rect 124462 99770 124490 100028
rect 123634 99742 123708 99770
rect 123576 99544 123628 99550
rect 123576 99486 123628 99492
rect 123588 96694 123616 99486
rect 123576 96688 123628 96694
rect 123576 96630 123628 96636
rect 123496 95118 123616 95146
rect 123484 94988 123536 94994
rect 123484 94930 123536 94936
rect 123312 94450 123432 94466
rect 123300 94444 123432 94450
rect 123352 94438 123432 94444
rect 123300 94386 123352 94392
rect 123392 94376 123444 94382
rect 123392 94318 123444 94324
rect 123300 94308 123352 94314
rect 123300 94250 123352 94256
rect 123312 21690 123340 94250
rect 123404 80714 123432 94318
rect 123496 82142 123524 94930
rect 123588 87854 123616 95118
rect 123576 87848 123628 87854
rect 123576 87790 123628 87796
rect 123680 87786 123708 99742
rect 123772 99742 123846 99770
rect 124416 99754 124490 99770
rect 124036 99748 124088 99754
rect 123772 94246 123800 99742
rect 124036 99690 124088 99696
rect 124312 99748 124364 99754
rect 124312 99690 124364 99696
rect 124404 99748 124490 99754
rect 124456 99742 124490 99748
rect 124554 99770 124582 100028
rect 124646 99929 124674 100028
rect 124738 100026 124766 100028
rect 124726 100020 124778 100026
rect 124726 99962 124778 99968
rect 124632 99920 124688 99929
rect 124830 99906 124858 100028
rect 124632 99855 124688 99864
rect 124784 99878 124858 99906
rect 124680 99816 124732 99822
rect 124554 99742 124628 99770
rect 124680 99758 124732 99764
rect 124404 99690 124456 99696
rect 123852 99680 123904 99686
rect 123852 99622 123904 99628
rect 123944 99680 123996 99686
rect 123944 99622 123996 99628
rect 123864 96082 123892 99622
rect 123956 97617 123984 99622
rect 124048 98297 124076 99690
rect 124220 99544 124272 99550
rect 124220 99486 124272 99492
rect 124034 98288 124090 98297
rect 124034 98223 124090 98232
rect 123942 97608 123998 97617
rect 123942 97543 123998 97552
rect 123852 96076 123904 96082
rect 123852 96018 123904 96024
rect 123760 94240 123812 94246
rect 123760 94182 123812 94188
rect 123668 87780 123720 87786
rect 123668 87722 123720 87728
rect 123484 82136 123536 82142
rect 123484 82078 123536 82084
rect 123392 80708 123444 80714
rect 123392 80650 123444 80656
rect 123300 21684 123352 21690
rect 123300 21626 123352 21632
rect 123208 21616 123260 21622
rect 123208 21558 123260 21564
rect 123116 21548 123168 21554
rect 123116 21490 123168 21496
rect 123024 18692 123076 18698
rect 123024 18634 123076 18640
rect 122932 6384 122984 6390
rect 122932 6326 122984 6332
rect 122840 5024 122892 5030
rect 122840 4966 122892 4972
rect 124232 4894 124260 99486
rect 124324 4962 124352 99690
rect 124496 99680 124548 99686
rect 124402 99648 124458 99657
rect 124496 99622 124548 99628
rect 124402 99583 124458 99592
rect 124416 94314 124444 99583
rect 124508 97306 124536 99622
rect 124496 97300 124548 97306
rect 124496 97242 124548 97248
rect 124496 94444 124548 94450
rect 124496 94386 124548 94392
rect 124404 94308 124456 94314
rect 124404 94250 124456 94256
rect 124404 94172 124456 94178
rect 124404 94114 124456 94120
rect 124416 7614 124444 94114
rect 124508 7682 124536 94386
rect 124600 7750 124628 99742
rect 124692 18630 124720 99758
rect 124784 94450 124812 99878
rect 124922 99804 124950 100028
rect 124876 99776 124950 99804
rect 124772 94444 124824 94450
rect 124772 94386 124824 94392
rect 124772 94308 124824 94314
rect 124772 94250 124824 94256
rect 124784 21486 124812 94250
rect 124876 35222 124904 99776
rect 125014 99668 125042 100028
rect 124968 99640 125042 99668
rect 124968 39438 124996 99640
rect 125106 99600 125134 100028
rect 125198 99770 125226 100028
rect 125290 99929 125318 100028
rect 125276 99920 125332 99929
rect 125276 99855 125332 99864
rect 125382 99770 125410 100028
rect 125198 99742 125272 99770
rect 125060 99572 125134 99600
rect 125060 94178 125088 99572
rect 125244 96801 125272 99742
rect 125336 99742 125410 99770
rect 125230 96792 125286 96801
rect 125230 96727 125286 96736
rect 125140 96688 125192 96694
rect 125336 96665 125364 99742
rect 125474 99668 125502 100028
rect 125566 99958 125594 100028
rect 125658 99963 125686 100028
rect 125554 99952 125606 99958
rect 125554 99894 125606 99900
rect 125644 99954 125700 99963
rect 125644 99889 125700 99898
rect 125842 99822 125870 100028
rect 125934 99963 125962 100028
rect 125920 99954 125976 99963
rect 126026 99958 126054 100028
rect 125920 99889 125976 99898
rect 126014 99952 126066 99958
rect 126014 99894 126066 99900
rect 125830 99816 125882 99822
rect 125830 99758 125882 99764
rect 125428 99640 125502 99668
rect 126118 99668 126146 100028
rect 126210 99963 126238 100028
rect 126196 99954 126252 99963
rect 126302 99958 126330 100028
rect 126394 99958 126422 100028
rect 126486 99963 126514 100028
rect 126196 99889 126252 99898
rect 126290 99952 126342 99958
rect 126290 99894 126342 99900
rect 126382 99952 126434 99958
rect 126382 99894 126434 99900
rect 126472 99954 126528 99963
rect 126472 99889 126528 99898
rect 126244 99748 126296 99754
rect 126244 99690 126296 99696
rect 125874 99648 125930 99657
rect 125428 97073 125456 99640
rect 126118 99640 126192 99668
rect 126256 99657 126284 99690
rect 126578 99668 126606 100028
rect 126670 99963 126698 100028
rect 126656 99954 126712 99963
rect 126656 99889 126712 99898
rect 126762 99668 126790 100028
rect 126854 99890 126882 100028
rect 126946 99958 126974 100028
rect 127038 99958 127066 100028
rect 127222 99958 127250 100028
rect 126934 99952 126986 99958
rect 126934 99894 126986 99900
rect 127026 99952 127078 99958
rect 127026 99894 127078 99900
rect 127210 99952 127262 99958
rect 127210 99894 127262 99900
rect 126842 99884 126894 99890
rect 126842 99826 126894 99832
rect 127072 99748 127124 99754
rect 127314 99736 127342 100028
rect 127420 100014 127572 100042
rect 127808 100030 127860 100036
rect 127314 99708 127388 99736
rect 127072 99690 127124 99696
rect 125874 99583 125930 99592
rect 125968 99612 126020 99618
rect 125506 99512 125562 99521
rect 125506 99447 125562 99456
rect 125782 99512 125838 99521
rect 125782 99447 125838 99456
rect 125414 97064 125470 97073
rect 125414 96999 125470 97008
rect 125140 96630 125192 96636
rect 125322 96656 125378 96665
rect 125048 94172 125100 94178
rect 125048 94114 125100 94120
rect 125046 92440 125102 92449
rect 125046 92375 125102 92384
rect 125060 92206 125088 92375
rect 125048 92200 125100 92206
rect 125048 92142 125100 92148
rect 125060 91118 125088 92142
rect 125152 91798 125180 96630
rect 125322 96591 125378 96600
rect 125520 96014 125548 99447
rect 125692 99408 125744 99414
rect 125598 99376 125654 99385
rect 125692 99350 125744 99356
rect 125598 99311 125654 99320
rect 125508 96008 125560 96014
rect 125508 95950 125560 95956
rect 125140 91792 125192 91798
rect 125140 91734 125192 91740
rect 125048 91112 125100 91118
rect 125048 91054 125100 91060
rect 124956 39432 125008 39438
rect 124956 39374 125008 39380
rect 124864 35216 124916 35222
rect 124864 35158 124916 35164
rect 124772 21480 124824 21486
rect 124772 21422 124824 21428
rect 124680 18624 124732 18630
rect 124680 18566 124732 18572
rect 124588 7744 124640 7750
rect 124588 7686 124640 7692
rect 124496 7676 124548 7682
rect 124496 7618 124548 7624
rect 124404 7608 124456 7614
rect 124404 7550 124456 7556
rect 124312 4956 124364 4962
rect 124312 4898 124364 4904
rect 124220 4888 124272 4894
rect 124220 4830 124272 4836
rect 125612 4826 125640 99311
rect 125704 6322 125732 99350
rect 125796 10334 125824 99447
rect 125888 11762 125916 99583
rect 125968 99554 126020 99560
rect 125980 15978 126008 99554
rect 126164 99414 126192 99640
rect 126242 99648 126298 99657
rect 126578 99640 126652 99668
rect 126242 99583 126298 99592
rect 126428 99612 126480 99618
rect 126428 99554 126480 99560
rect 126244 99544 126296 99550
rect 126440 99498 126468 99554
rect 126244 99486 126296 99492
rect 126152 99408 126204 99414
rect 126152 99350 126204 99356
rect 126150 99240 126206 99249
rect 126150 99175 126206 99184
rect 126058 98288 126114 98297
rect 126058 98223 126114 98232
rect 126072 20126 126100 98223
rect 126164 21418 126192 99175
rect 126256 39370 126284 99486
rect 126348 99470 126468 99498
rect 126520 99544 126572 99550
rect 126520 99486 126572 99492
rect 126348 87650 126376 99470
rect 126428 99408 126480 99414
rect 126428 99350 126480 99356
rect 126440 87718 126468 99350
rect 126532 95946 126560 99486
rect 126624 97345 126652 99640
rect 126716 99640 126790 99668
rect 126716 98161 126744 99640
rect 126888 99612 126940 99618
rect 126888 99554 126940 99560
rect 126900 98297 126928 99554
rect 126886 98288 126942 98297
rect 126886 98223 126942 98232
rect 126702 98152 126758 98161
rect 126702 98087 126758 98096
rect 127084 97510 127112 99690
rect 127256 99612 127308 99618
rect 127256 99554 127308 99560
rect 127072 97504 127124 97510
rect 127072 97446 127124 97452
rect 126610 97336 126666 97345
rect 126610 97271 126666 97280
rect 126520 95940 126572 95946
rect 126520 95882 126572 95888
rect 126980 95056 127032 95062
rect 126980 94998 127032 95004
rect 126428 87712 126480 87718
rect 126428 87654 126480 87660
rect 126336 87644 126388 87650
rect 126336 87586 126388 87592
rect 126244 39364 126296 39370
rect 126244 39306 126296 39312
rect 126152 21412 126204 21418
rect 126152 21354 126204 21360
rect 126060 20120 126112 20126
rect 126060 20062 126112 20068
rect 126992 16574 127020 94998
rect 127268 88942 127296 99554
rect 127360 98326 127388 99708
rect 127348 98320 127400 98326
rect 127348 98262 127400 98268
rect 127544 89714 127572 100014
rect 127624 99884 127676 99890
rect 127624 99826 127676 99832
rect 127452 89686 127572 89714
rect 127256 88936 127308 88942
rect 127256 88878 127308 88884
rect 127452 19990 127480 89686
rect 127532 88936 127584 88942
rect 127532 88878 127584 88884
rect 127440 19984 127492 19990
rect 127440 19926 127492 19932
rect 126992 16546 127480 16574
rect 125968 15972 126020 15978
rect 125968 15914 126020 15920
rect 125876 11756 125928 11762
rect 125876 11698 125928 11704
rect 125784 10328 125836 10334
rect 125784 10270 125836 10276
rect 125692 6316 125744 6322
rect 125692 6258 125744 6264
rect 125600 4820 125652 4826
rect 125600 4762 125652 4768
rect 126888 3800 126940 3806
rect 126888 3742 126940 3748
rect 123576 3732 123628 3738
rect 123576 3674 123628 3680
rect 122564 3528 122616 3534
rect 122564 3470 122616 3476
rect 123588 480 123616 3674
rect 125784 3664 125836 3670
rect 125784 3606 125836 3612
rect 124678 3360 124734 3369
rect 124678 3295 124734 3304
rect 124692 480 124720 3295
rect 125796 480 125824 3606
rect 126900 480 126928 3742
rect 127452 3482 127480 16546
rect 127544 6186 127572 88878
rect 127636 6254 127664 99826
rect 127716 98320 127768 98326
rect 127716 98262 127768 98268
rect 127728 15910 127756 98262
rect 127820 20058 127848 100030
rect 128096 99346 128124 149534
rect 128188 100366 128216 151778
rect 128176 100360 128228 100366
rect 128176 100302 128228 100308
rect 128084 99340 128136 99346
rect 128084 99282 128136 99288
rect 127992 96756 128044 96762
rect 127992 96698 128044 96704
rect 127900 96552 127952 96558
rect 127900 96494 127952 96500
rect 127808 20052 127860 20058
rect 127808 19994 127860 20000
rect 127716 15904 127768 15910
rect 127716 15846 127768 15852
rect 127624 6248 127676 6254
rect 127624 6190 127676 6196
rect 127532 6180 127584 6186
rect 127532 6122 127584 6128
rect 127912 3806 127940 96494
rect 127900 3800 127952 3806
rect 127900 3742 127952 3748
rect 128004 3670 128032 96698
rect 128084 93832 128136 93838
rect 128084 93774 128136 93780
rect 128096 3738 128124 93774
rect 128372 89842 128400 152050
rect 128280 89814 128400 89842
rect 128280 89298 128308 89814
rect 128360 89684 128412 89690
rect 128360 89626 128412 89632
rect 128372 89418 128400 89626
rect 128360 89412 128412 89418
rect 128360 89354 128412 89360
rect 128280 89270 128400 89298
rect 128372 85542 128400 89270
rect 128464 88330 128492 152118
rect 128452 88324 128504 88330
rect 128452 88266 128504 88272
rect 128556 88262 128584 152186
rect 128636 151904 128688 151910
rect 128636 151846 128688 151852
rect 128648 89418 128676 151846
rect 128740 91050 128768 152866
rect 136086 152552 136142 152561
rect 136086 152487 136142 152496
rect 128820 152040 128872 152046
rect 128820 151982 128872 151988
rect 128832 92478 128860 151982
rect 128912 151972 128964 151978
rect 128912 151914 128964 151920
rect 128820 92472 128872 92478
rect 128820 92414 128872 92420
rect 128832 92206 128860 92414
rect 128820 92200 128872 92206
rect 128820 92142 128872 92148
rect 128924 92138 128952 151914
rect 129830 151872 129886 151881
rect 129830 151807 129886 151816
rect 129004 150816 129056 150822
rect 129004 150758 129056 150764
rect 129016 133890 129044 150758
rect 129004 133884 129056 133890
rect 129004 133826 129056 133832
rect 129188 97980 129240 97986
rect 129188 97922 129240 97928
rect 129096 97232 129148 97238
rect 129096 97174 129148 97180
rect 129004 96620 129056 96626
rect 129004 96562 129056 96568
rect 128912 92132 128964 92138
rect 128912 92074 128964 92080
rect 128728 91044 128780 91050
rect 128728 90986 128780 90992
rect 128740 90642 128768 90986
rect 128728 90636 128780 90642
rect 128728 90578 128780 90584
rect 128636 89412 128688 89418
rect 128636 89354 128688 89360
rect 128544 88256 128596 88262
rect 128544 88198 128596 88204
rect 128360 85536 128412 85542
rect 128360 85478 128412 85484
rect 129016 3874 129044 96562
rect 129108 53106 129136 97174
rect 129200 53174 129228 97922
rect 129740 97912 129792 97918
rect 129740 97854 129792 97860
rect 129280 97164 129332 97170
rect 129280 97106 129332 97112
rect 129292 54534 129320 97106
rect 129280 54528 129332 54534
rect 129280 54470 129332 54476
rect 129188 53168 129240 53174
rect 129188 53110 129240 53116
rect 129096 53100 129148 53106
rect 129096 53042 129148 53048
rect 129752 16574 129780 97854
rect 129844 89350 129872 151807
rect 131120 97844 131172 97850
rect 131120 97786 131172 97792
rect 129832 89344 129884 89350
rect 129832 89286 129884 89292
rect 129752 16546 130240 16574
rect 129096 6588 129148 6594
rect 129096 6530 129148 6536
rect 129004 3868 129056 3874
rect 129004 3810 129056 3816
rect 128084 3732 128136 3738
rect 128084 3674 128136 3680
rect 127992 3664 128044 3670
rect 127992 3606 128044 3612
rect 127452 3454 128032 3482
rect 128004 480 128032 3454
rect 129108 480 129136 6530
rect 130212 480 130240 16546
rect 131132 3482 131160 97786
rect 131764 97776 131816 97782
rect 131764 97718 131816 97724
rect 131212 42152 131264 42158
rect 131212 42094 131264 42100
rect 131224 4146 131252 42094
rect 131212 4140 131264 4146
rect 131212 4082 131264 4088
rect 131132 3454 131344 3482
rect 131316 480 131344 3454
rect 131776 3262 131804 97718
rect 133880 97708 133932 97714
rect 133880 97650 133932 97656
rect 133892 16574 133920 97650
rect 135904 97640 135956 97646
rect 135904 97582 135956 97588
rect 133892 16546 134656 16574
rect 132408 4140 132460 4146
rect 132408 4082 132460 4088
rect 131764 3256 131816 3262
rect 131764 3198 131816 3204
rect 132420 480 132448 4082
rect 133512 3256 133564 3262
rect 133512 3198 133564 3204
rect 133524 480 133552 3198
rect 134628 480 134656 16546
rect 135720 3936 135772 3942
rect 135720 3878 135772 3884
rect 135732 480 135760 3878
rect 135916 3398 135944 97582
rect 135996 96416 136048 96422
rect 135996 96358 136048 96364
rect 136008 3942 136036 96358
rect 136100 71738 136128 152487
rect 138662 152416 138718 152425
rect 138662 152351 138718 152360
rect 138676 118658 138704 152351
rect 580356 151088 580408 151094
rect 580356 151030 580408 151036
rect 580172 150476 580224 150482
rect 580172 150418 580224 150424
rect 580184 148617 580212 150418
rect 580264 149456 580316 149462
rect 580264 149398 580316 149404
rect 580170 148608 580226 148617
rect 580170 148543 580226 148552
rect 579988 133884 580040 133890
rect 579988 133826 580040 133832
rect 580000 132977 580028 133826
rect 579986 132968 580042 132977
rect 579986 132903 580042 132912
rect 138664 118652 138716 118658
rect 138664 118594 138716 118600
rect 580172 118652 580224 118658
rect 580172 118594 580224 118600
rect 580184 117337 580212 118594
rect 580170 117328 580226 117337
rect 580170 117263 580226 117272
rect 200764 97572 200816 97578
rect 200764 97514 200816 97520
rect 176660 96348 176712 96354
rect 176660 96290 176712 96296
rect 162124 94920 162176 94926
rect 162124 94862 162176 94868
rect 153198 94752 153254 94761
rect 153198 94687 153254 94696
rect 142160 92404 142212 92410
rect 142160 92346 142212 92352
rect 136088 71732 136140 71738
rect 136088 71674 136140 71680
rect 136732 42084 136784 42090
rect 136732 42026 136784 42032
rect 136744 16574 136772 42026
rect 140778 40896 140834 40905
rect 140778 40831 140834 40840
rect 139398 19000 139454 19009
rect 139398 18935 139454 18944
rect 139412 16574 139440 18935
rect 140792 16574 140820 40831
rect 136744 16546 136864 16574
rect 139412 16546 140176 16574
rect 140792 16546 141280 16574
rect 135996 3936 136048 3942
rect 135996 3878 136048 3884
rect 135904 3392 135956 3398
rect 135904 3334 135956 3340
rect 136836 480 136864 16546
rect 139032 4004 139084 4010
rect 139032 3946 139084 3952
rect 137928 3392 137980 3398
rect 137928 3334 137980 3340
rect 137940 480 137968 3334
rect 139044 480 139072 3946
rect 140148 480 140176 16546
rect 141252 480 141280 16546
rect 142172 3482 142200 92346
rect 144920 89616 144972 89622
rect 144920 89558 144972 89564
rect 142252 24540 142304 24546
rect 142252 24482 142304 24488
rect 142264 4010 142292 24482
rect 143540 17672 143592 17678
rect 143540 17614 143592 17620
rect 143552 16574 143580 17614
rect 144932 16574 144960 89558
rect 149060 27328 149112 27334
rect 149060 27270 149112 27276
rect 146300 26104 146352 26110
rect 146300 26046 146352 26052
rect 146312 16574 146340 26046
rect 147680 21888 147732 21894
rect 147680 21830 147732 21836
rect 143552 16546 144592 16574
rect 144932 16546 145696 16574
rect 146312 16546 146800 16574
rect 142252 4004 142304 4010
rect 142252 3946 142304 3952
rect 143448 4004 143500 4010
rect 143448 3946 143500 3952
rect 142172 3454 142384 3482
rect 142356 480 142384 3454
rect 143460 480 143488 3946
rect 144564 480 144592 16546
rect 145668 480 145696 16546
rect 146772 480 146800 16546
rect 147692 3482 147720 21830
rect 149072 16574 149100 27270
rect 150440 27260 150492 27266
rect 150440 27202 150492 27208
rect 150452 16574 150480 27202
rect 149072 16546 150112 16574
rect 150452 16546 151216 16574
rect 147772 10804 147824 10810
rect 147772 10746 147824 10752
rect 147784 4010 147812 10746
rect 147772 4004 147824 4010
rect 147772 3946 147824 3952
rect 148968 4004 149020 4010
rect 148968 3946 149020 3952
rect 147692 3454 147904 3482
rect 147876 480 147904 3454
rect 148980 480 149008 3946
rect 150084 480 150112 16546
rect 151188 480 151216 16546
rect 152280 12232 152332 12238
rect 152280 12174 152332 12180
rect 152292 480 152320 12174
rect 153212 3398 153240 94687
rect 158720 90704 158772 90710
rect 158720 90646 158772 90652
rect 157338 42120 157394 42129
rect 157338 42055 157394 42064
rect 153290 28520 153346 28529
rect 153290 28455 153346 28464
rect 153304 16574 153332 28455
rect 157352 16574 157380 42055
rect 153304 16546 153424 16574
rect 157352 16546 157840 16574
rect 153200 3392 153252 3398
rect 153200 3334 153252 3340
rect 153396 480 153424 16546
rect 155592 13524 155644 13530
rect 155592 13466 155644 13472
rect 154488 3392 154540 3398
rect 154488 3334 154540 3340
rect 154500 480 154528 3334
rect 155604 480 155632 13466
rect 156694 11792 156750 11801
rect 156694 11727 156750 11736
rect 156708 480 156736 11727
rect 157812 480 157840 16546
rect 158732 3482 158760 90646
rect 158812 31544 158864 31550
rect 158812 31486 158864 31492
rect 158824 4010 158852 31486
rect 160100 30184 160152 30190
rect 160100 30126 160152 30132
rect 160112 16574 160140 30126
rect 160112 16546 161152 16574
rect 158812 4004 158864 4010
rect 158812 3946 158864 3952
rect 160008 4004 160060 4010
rect 160008 3946 160060 3952
rect 158732 3454 158944 3482
rect 158916 480 158944 3454
rect 160020 480 160048 3946
rect 161124 480 161152 16546
rect 162032 16312 162084 16318
rect 162032 16254 162084 16260
rect 162044 3482 162072 16254
rect 162136 4146 162164 94862
rect 171140 92336 171192 92342
rect 171140 92278 171192 92284
rect 164240 85196 164292 85202
rect 164240 85138 164292 85144
rect 162860 31476 162912 31482
rect 162860 31418 162912 31424
rect 162872 16574 162900 31418
rect 162872 16546 163360 16574
rect 162124 4140 162176 4146
rect 162124 4082 162176 4088
rect 162044 3454 162256 3482
rect 162228 480 162256 3454
rect 163332 480 163360 16546
rect 164148 3868 164200 3874
rect 164148 3810 164200 3816
rect 164160 3398 164188 3810
rect 164252 3482 164280 85138
rect 165620 41200 165672 41206
rect 165620 41142 165672 41148
rect 164332 17604 164384 17610
rect 164332 17546 164384 17552
rect 164344 3874 164372 17546
rect 165632 16574 165660 41142
rect 169850 40760 169906 40769
rect 169850 40695 169906 40704
rect 169024 19032 169076 19038
rect 169024 18974 169076 18980
rect 168380 18964 168432 18970
rect 168380 18906 168432 18912
rect 168392 16574 168420 18906
rect 165632 16546 166672 16574
rect 168392 16546 168880 16574
rect 164332 3868 164384 3874
rect 164332 3810 164384 3816
rect 165528 3868 165580 3874
rect 165528 3810 165580 3816
rect 164252 3454 164464 3482
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 164436 480 164464 3454
rect 165540 480 165568 3810
rect 166644 480 166672 16546
rect 167736 3392 167788 3398
rect 167736 3334 167788 3340
rect 167748 480 167776 3334
rect 168852 480 168880 16546
rect 169036 3874 169064 18974
rect 169864 16574 169892 40695
rect 171152 16574 171180 92278
rect 175280 92268 175332 92274
rect 175280 92210 175332 92216
rect 173898 36408 173954 36417
rect 173898 36343 173954 36352
rect 172518 20088 172574 20097
rect 172518 20023 172574 20032
rect 172532 16574 172560 20023
rect 173912 16574 173940 36343
rect 169864 16546 169984 16574
rect 171152 16546 172192 16574
rect 172532 16546 173296 16574
rect 173912 16546 174400 16574
rect 169024 3868 169076 3874
rect 169024 3810 169076 3816
rect 169956 480 169984 16546
rect 170956 4072 171008 4078
rect 170956 4014 171008 4020
rect 170968 2122 170996 4014
rect 170968 2094 171088 2122
rect 171060 480 171088 2094
rect 172164 480 172192 16546
rect 173268 480 173296 16546
rect 174372 480 174400 16546
rect 175292 3482 175320 92210
rect 175372 21820 175424 21826
rect 175372 21762 175424 21768
rect 175384 4078 175412 21762
rect 176672 16574 176700 96290
rect 193220 96280 193272 96286
rect 193220 96222 193272 96228
rect 191840 91112 191892 91118
rect 191840 91054 191892 91060
rect 178040 89548 178092 89554
rect 178040 89490 178092 89496
rect 178052 16574 178080 89490
rect 180800 89480 180852 89486
rect 180800 89422 180852 89428
rect 179420 23180 179472 23186
rect 179420 23122 179472 23128
rect 179432 16574 179460 23122
rect 176672 16546 177712 16574
rect 178052 16546 178816 16574
rect 179432 16546 179920 16574
rect 175372 4072 175424 4078
rect 175372 4014 175424 4020
rect 176568 4072 176620 4078
rect 176568 4014 176620 4020
rect 175292 3454 175504 3482
rect 175476 480 175504 3454
rect 176580 480 176608 4014
rect 177684 480 177712 16546
rect 178788 480 178816 16546
rect 179892 480 179920 16546
rect 180812 3398 180840 89422
rect 190458 40624 190514 40633
rect 190458 40559 190514 40568
rect 186318 37224 186374 37233
rect 186318 37159 186374 37168
rect 180892 36712 180944 36718
rect 180892 36654 180944 36660
rect 180904 16574 180932 36654
rect 182180 23112 182232 23118
rect 182180 23054 182232 23060
rect 182192 16574 182220 23054
rect 183560 18896 183612 18902
rect 183560 18838 183612 18844
rect 183572 16574 183600 18838
rect 180904 16546 181024 16574
rect 182192 16546 183232 16574
rect 183572 16546 184336 16574
rect 180800 3392 180852 3398
rect 180800 3334 180852 3340
rect 180996 480 181024 16546
rect 182088 3392 182140 3398
rect 182088 3334 182140 3340
rect 182100 480 182128 3334
rect 183204 480 183232 16546
rect 184308 480 184336 16546
rect 185400 6520 185452 6526
rect 185400 6462 185452 6468
rect 185412 480 185440 6462
rect 186332 3398 186360 37159
rect 190472 16574 190500 40559
rect 190472 16546 190960 16574
rect 189814 7576 189870 7585
rect 189814 7511 189870 7520
rect 188712 6452 188764 6458
rect 188712 6394 188764 6400
rect 186504 5364 186556 5370
rect 186504 5306 186556 5312
rect 186320 3392 186372 3398
rect 186320 3334 186372 3340
rect 186516 480 186544 5306
rect 187608 3392 187660 3398
rect 187608 3334 187660 3340
rect 187620 480 187648 3334
rect 188724 480 188752 6394
rect 189828 480 189856 7511
rect 190932 480 190960 16546
rect 191852 3482 191880 91054
rect 191932 23044 191984 23050
rect 191932 22986 191984 22992
rect 191944 4078 191972 22986
rect 193232 16574 193260 96222
rect 200120 96212 200172 96218
rect 200120 96154 200172 96160
rect 194600 92200 194652 92206
rect 194600 92142 194652 92148
rect 194612 16574 194640 92142
rect 197360 85264 197412 85270
rect 197360 85206 197412 85212
rect 195980 22976 196032 22982
rect 195980 22918 196032 22924
rect 195992 16574 196020 22918
rect 193232 16546 194272 16574
rect 194612 16546 195376 16574
rect 195992 16546 196480 16574
rect 191932 4072 191984 4078
rect 191932 4014 191984 4020
rect 193128 4072 193180 4078
rect 193128 4014 193180 4020
rect 191852 3454 192064 3482
rect 192036 480 192064 3454
rect 193140 480 193168 4014
rect 194244 480 194272 16546
rect 195348 480 195376 16546
rect 196452 480 196480 16546
rect 197372 3398 197400 85206
rect 197452 36644 197504 36650
rect 197452 36586 197504 36592
rect 197464 16574 197492 36586
rect 198740 24472 198792 24478
rect 198740 24414 198792 24420
rect 198752 16574 198780 24414
rect 200132 16574 200160 96154
rect 200776 88058 200804 97514
rect 209044 97504 209096 97510
rect 209044 97446 209096 97452
rect 208400 88324 208452 88330
rect 208400 88266 208452 88272
rect 200764 88052 200816 88058
rect 200764 87994 200816 88000
rect 207018 38312 207074 38321
rect 207018 38247 207074 38256
rect 202878 37088 202934 37097
rect 202878 37023 202934 37032
rect 197464 16546 197584 16574
rect 198752 16546 199792 16574
rect 200132 16546 200896 16574
rect 197360 3392 197412 3398
rect 197360 3334 197412 3340
rect 197556 480 197584 16546
rect 198648 3392 198700 3398
rect 198648 3334 198700 3340
rect 198660 480 198688 3334
rect 199764 480 199792 16546
rect 200868 480 200896 16546
rect 201960 8152 202012 8158
rect 201960 8094 202012 8100
rect 201972 480 202000 8094
rect 202892 3398 202920 37023
rect 207032 16574 207060 38247
rect 207032 16546 207520 16574
rect 203062 9480 203118 9489
rect 203062 9415 203118 9424
rect 202880 3392 202932 3398
rect 202880 3334 202932 3340
rect 203076 480 203104 9415
rect 206374 9344 206430 9353
rect 206374 9279 206430 9288
rect 205272 8084 205324 8090
rect 205272 8026 205324 8032
rect 204168 3392 204220 3398
rect 204168 3334 204220 3340
rect 204180 480 204208 3334
rect 205284 480 205312 8026
rect 206388 480 206416 9279
rect 207492 480 207520 16546
rect 208412 3482 208440 88266
rect 208492 24404 208544 24410
rect 208492 24346 208544 24352
rect 208504 4078 208532 24346
rect 209056 8974 209084 97446
rect 278044 97436 278096 97442
rect 278044 97378 278096 97384
rect 247040 94852 247092 94858
rect 247040 94794 247092 94800
rect 235998 94616 236054 94625
rect 235998 94551 236054 94560
rect 224960 92132 225012 92138
rect 224960 92074 225012 92080
rect 211160 90636 211212 90642
rect 211160 90578 211212 90584
rect 211172 16574 211200 90578
rect 218060 89412 218112 89418
rect 218060 89354 218112 89360
rect 216680 32904 216732 32910
rect 216680 32846 216732 32852
rect 212540 24336 212592 24342
rect 212540 24278 212592 24284
rect 212552 16574 212580 24278
rect 215300 24268 215352 24274
rect 215300 24210 215352 24216
rect 213920 20460 213972 20466
rect 213920 20402 213972 20408
rect 213932 16574 213960 20402
rect 215312 16574 215340 24210
rect 216692 16574 216720 32846
rect 218072 16574 218100 89354
rect 223578 38176 223634 38185
rect 223578 38111 223634 38120
rect 219438 24440 219494 24449
rect 219438 24375 219494 24384
rect 211172 16546 211936 16574
rect 212552 16546 213040 16574
rect 213932 16546 214144 16574
rect 215312 16546 216352 16574
rect 216692 16546 217456 16574
rect 218072 16546 218560 16574
rect 209044 8968 209096 8974
rect 209044 8910 209096 8916
rect 208492 4072 208544 4078
rect 208492 4014 208544 4020
rect 209688 4072 209740 4078
rect 209688 4014 209740 4020
rect 208412 3454 208624 3482
rect 208596 480 208624 3454
rect 209700 480 209728 4014
rect 210792 3936 210844 3942
rect 210792 3878 210844 3884
rect 210804 480 210832 3878
rect 211908 480 211936 16546
rect 213012 480 213040 16546
rect 214116 480 214144 16546
rect 215208 8016 215260 8022
rect 215208 7958 215260 7964
rect 215220 480 215248 7958
rect 216324 480 216352 16546
rect 217428 480 217456 16546
rect 218532 480 218560 16546
rect 219452 3482 219480 24375
rect 219530 21448 219586 21457
rect 219530 21383 219586 21392
rect 219544 3942 219572 21383
rect 223592 16574 223620 38111
rect 223592 16546 224080 16574
rect 221832 7948 221884 7954
rect 221832 7890 221884 7896
rect 219532 3936 219584 3942
rect 219532 3878 219584 3884
rect 220728 3936 220780 3942
rect 220728 3878 220780 3884
rect 219452 3454 219664 3482
rect 219636 480 219664 3454
rect 220740 480 220768 3878
rect 221844 480 221872 7890
rect 222934 6624 222990 6633
rect 222934 6559 222990 6568
rect 222948 480 222976 6559
rect 224052 480 224080 16546
rect 224972 3482 225000 92074
rect 227720 88256 227772 88262
rect 227720 88198 227772 88204
rect 225052 46232 225104 46238
rect 225052 46174 225104 46180
rect 225064 3942 225092 46174
rect 226340 21752 226392 21758
rect 226340 21694 226392 21700
rect 226352 16574 226380 21694
rect 227732 16574 227760 88198
rect 230480 38276 230532 38282
rect 230480 38218 230532 38224
rect 230492 16574 230520 38218
rect 233240 38208 233292 38214
rect 233240 38150 233292 38156
rect 233252 16574 233280 38150
rect 226352 16546 227392 16574
rect 227732 16546 228496 16574
rect 230492 16546 230704 16574
rect 233252 16546 234016 16574
rect 225052 3936 225104 3942
rect 225052 3878 225104 3884
rect 226248 3936 226300 3942
rect 226248 3878 226300 3884
rect 224972 3454 225184 3482
rect 225156 480 225184 3454
rect 226260 480 226288 3878
rect 227364 480 227392 16546
rect 228468 480 228496 16546
rect 229560 7880 229612 7886
rect 229560 7822 229612 7828
rect 229572 480 229600 7822
rect 230676 480 230704 16546
rect 231768 7812 231820 7818
rect 231768 7754 231820 7760
rect 231780 480 231808 7754
rect 232872 5296 232924 5302
rect 232872 5238 232924 5244
rect 232884 480 232912 5238
rect 233988 480 234016 16546
rect 235080 9308 235132 9314
rect 235080 9250 235132 9256
rect 235092 480 235120 9250
rect 236012 3398 236040 94551
rect 241520 89344 241572 89350
rect 241520 89286 241572 89292
rect 237380 39772 237432 39778
rect 237380 39714 237432 39720
rect 237392 16574 237420 39714
rect 240138 27160 240194 27169
rect 240138 27095 240194 27104
rect 240152 16574 240180 27095
rect 237392 16546 238432 16574
rect 240152 16546 240640 16574
rect 236182 9208 236238 9217
rect 236182 9143 236238 9152
rect 236000 3392 236052 3398
rect 236000 3334 236052 3340
rect 236196 480 236224 9143
rect 237288 3392 237340 3398
rect 237288 3334 237340 3340
rect 237300 480 237328 3334
rect 238404 480 238432 16546
rect 239494 9072 239550 9081
rect 239494 9007 239550 9016
rect 239508 480 239536 9007
rect 240612 480 240640 16546
rect 241532 3482 241560 89286
rect 244280 86624 244332 86630
rect 244280 86566 244332 86572
rect 242900 41132 242952 41138
rect 242900 41074 242952 41080
rect 241612 26036 241664 26042
rect 241612 25978 241664 25984
rect 241624 3942 241652 25978
rect 242912 16574 242940 41074
rect 244292 16574 244320 86566
rect 245660 25968 245712 25974
rect 245660 25910 245712 25916
rect 245672 16574 245700 25910
rect 242912 16546 243952 16574
rect 244292 16546 245056 16574
rect 245672 16546 246160 16574
rect 241612 3936 241664 3942
rect 241612 3878 241664 3884
rect 242808 3936 242860 3942
rect 242808 3878 242860 3884
rect 241532 3454 241744 3482
rect 241716 480 241744 3454
rect 242820 480 242848 3878
rect 243924 480 243952 16546
rect 245028 480 245056 16546
rect 246132 480 246160 16546
rect 247052 3482 247080 94794
rect 252560 94784 252612 94790
rect 252560 94726 252612 94732
rect 251180 88188 251232 88194
rect 251180 88130 251232 88136
rect 247132 86556 247184 86562
rect 247132 86498 247184 86504
rect 247144 3942 247172 86498
rect 248420 25900 248472 25906
rect 248420 25842 248472 25848
rect 248432 16574 248460 25842
rect 249800 22908 249852 22914
rect 249800 22850 249852 22856
rect 249812 16574 249840 22850
rect 251192 16574 251220 88130
rect 248432 16546 249472 16574
rect 249812 16546 250576 16574
rect 251192 16546 251680 16574
rect 247132 3936 247184 3942
rect 247132 3878 247184 3884
rect 248328 3936 248380 3942
rect 248328 3878 248380 3884
rect 247052 3454 247264 3482
rect 247236 480 247264 3454
rect 248340 480 248368 3878
rect 249444 480 249472 16546
rect 250548 480 250576 16546
rect 251652 480 251680 16546
rect 252572 3398 252600 94726
rect 266360 94716 266412 94722
rect 266360 94658 266412 94664
rect 258080 89276 258132 89282
rect 258080 89218 258132 89224
rect 252652 25832 252704 25838
rect 252652 25774 252704 25780
rect 252664 16574 252692 25774
rect 255318 25528 255374 25537
rect 255318 25463 255374 25472
rect 255332 16574 255360 25463
rect 256698 22944 256754 22953
rect 256698 22879 256754 22888
rect 256712 16574 256740 22879
rect 252664 16546 252784 16574
rect 255332 16546 256096 16574
rect 256712 16546 257200 16574
rect 252560 3392 252612 3398
rect 252560 3334 252612 3340
rect 252756 480 252784 16546
rect 254950 8936 255006 8945
rect 254950 8871 255006 8880
rect 253848 3392 253900 3398
rect 253848 3334 253900 3340
rect 253860 480 253888 3334
rect 254964 480 254992 8871
rect 256068 480 256096 16546
rect 257172 480 257200 16546
rect 258092 3482 258120 89218
rect 258172 27192 258224 27198
rect 258172 27134 258224 27140
rect 258184 3942 258212 27134
rect 262220 27124 262272 27130
rect 262220 27066 262272 27072
rect 259460 22840 259512 22846
rect 259460 22782 259512 22788
rect 259472 16574 259500 22782
rect 262232 16574 262260 27066
rect 264980 27056 265032 27062
rect 264980 26998 265032 27004
rect 263600 22772 263652 22778
rect 263600 22714 263652 22720
rect 263612 16574 263640 22714
rect 264992 16574 265020 26998
rect 266372 16574 266400 94658
rect 274640 86488 274692 86494
rect 274640 86430 274692 86436
rect 270498 84960 270554 84969
rect 270498 84895 270554 84904
rect 269118 27024 269174 27033
rect 269118 26959 269174 26968
rect 259472 16546 260512 16574
rect 262232 16546 262720 16574
rect 263612 16546 263824 16574
rect 264992 16546 266032 16574
rect 266372 16546 267136 16574
rect 258172 3936 258224 3942
rect 258172 3878 258224 3884
rect 259368 3936 259420 3942
rect 259368 3878 259420 3884
rect 258092 3454 258304 3482
rect 258276 480 258304 3454
rect 259380 480 259408 3878
rect 260484 480 260512 16546
rect 261576 9240 261628 9246
rect 261576 9182 261628 9188
rect 261588 480 261616 9182
rect 262692 480 262720 16546
rect 263796 480 263824 16546
rect 264888 9172 264940 9178
rect 264888 9114 264940 9120
rect 264900 480 264928 9114
rect 266004 480 266032 16546
rect 267108 480 267136 16546
rect 268200 9104 268252 9110
rect 268200 9046 268252 9052
rect 268212 480 268240 9046
rect 269132 3398 269160 26959
rect 270512 16574 270540 84895
rect 273258 26888 273314 26897
rect 273258 26823 273314 26832
rect 273272 16574 273300 26823
rect 270512 16546 271552 16574
rect 273272 16546 273760 16574
rect 269304 10736 269356 10742
rect 269304 10678 269356 10684
rect 269120 3392 269172 3398
rect 269120 3334 269172 3340
rect 269316 480 269344 10678
rect 270408 3392 270460 3398
rect 270408 3334 270460 3340
rect 270420 480 270448 3334
rect 271524 480 271552 16546
rect 272614 10432 272670 10441
rect 272614 10367 272670 10376
rect 272628 480 272656 10367
rect 273732 480 273760 16546
rect 274652 3482 274680 86430
rect 276020 28688 276072 28694
rect 276020 28630 276072 28636
rect 274732 26988 274784 26994
rect 274732 26930 274784 26936
rect 274744 3942 274772 26930
rect 276032 16574 276060 28630
rect 276032 16546 277072 16574
rect 274732 3936 274784 3942
rect 274732 3878 274784 3884
rect 275928 3936 275980 3942
rect 275928 3878 275980 3884
rect 274652 3454 274864 3482
rect 274836 480 274864 3454
rect 275940 480 275968 3878
rect 277044 480 277072 16546
rect 278056 4010 278084 97378
rect 295984 97368 296036 97374
rect 295984 97310 296036 97316
rect 289818 94480 289874 94489
rect 289818 94415 289874 94424
rect 287060 89208 287112 89214
rect 287060 89150 287112 89156
rect 282920 86420 282972 86426
rect 282920 86362 282972 86368
rect 280160 28620 280212 28626
rect 280160 28562 280212 28568
rect 278780 26920 278832 26926
rect 278780 26862 278832 26868
rect 278792 16574 278820 26862
rect 278792 16546 279280 16574
rect 278136 9036 278188 9042
rect 278136 8978 278188 8984
rect 278044 4004 278096 4010
rect 278044 3946 278096 3952
rect 278148 480 278176 8978
rect 279252 480 279280 16546
rect 280172 3482 280200 28562
rect 281540 28552 281592 28558
rect 281540 28494 281592 28500
rect 281552 16574 281580 28494
rect 282932 16574 282960 86362
rect 285770 28384 285826 28393
rect 285770 28319 285826 28328
rect 285678 28248 285734 28257
rect 285678 28183 285734 28192
rect 281552 16546 282592 16574
rect 282932 16546 283696 16574
rect 280252 10668 280304 10674
rect 280252 10610 280304 10616
rect 280264 3942 280292 10610
rect 280252 3936 280304 3942
rect 280252 3878 280304 3884
rect 281448 3936 281500 3942
rect 281448 3878 281500 3884
rect 280172 3454 280384 3482
rect 280356 480 280384 3454
rect 281460 480 281488 3878
rect 282564 480 282592 16546
rect 283668 480 283696 16546
rect 284760 10600 284812 10606
rect 284760 10542 284812 10548
rect 284772 480 284800 10542
rect 285692 3398 285720 28183
rect 285784 16574 285812 28319
rect 287072 16574 287100 89150
rect 289832 16574 289860 94415
rect 291200 90568 291252 90574
rect 291200 90510 291252 90516
rect 285784 16546 285904 16574
rect 287072 16546 288112 16574
rect 289832 16546 290320 16574
rect 285680 3392 285732 3398
rect 285680 3334 285732 3340
rect 285876 480 285904 16546
rect 286968 3392 287020 3398
rect 286968 3334 287020 3340
rect 286980 480 287008 3334
rect 288084 480 288112 16546
rect 289174 10296 289230 10305
rect 289174 10231 289230 10240
rect 289188 480 289216 10231
rect 290292 480 290320 16546
rect 291212 3482 291240 90510
rect 293960 89140 294012 89146
rect 293960 89082 294012 89088
rect 291292 28484 291344 28490
rect 291292 28426 291344 28432
rect 291304 4010 291332 28426
rect 293972 16574 294000 89082
rect 295340 28416 295392 28422
rect 295340 28358 295392 28364
rect 295352 16574 295380 28358
rect 293972 16546 294736 16574
rect 295352 16546 295840 16574
rect 293592 4072 293644 4078
rect 293592 4014 293644 4020
rect 291292 4004 291344 4010
rect 291292 3946 291344 3952
rect 292488 4004 292540 4010
rect 292488 3946 292540 3952
rect 291212 3454 291424 3482
rect 291396 480 291424 3454
rect 292500 480 292528 3946
rect 293604 480 293632 4014
rect 294708 480 294736 16546
rect 295812 480 295840 16546
rect 295996 4010 296024 97310
rect 446404 97300 446456 97306
rect 446404 97242 446456 97248
rect 296720 94648 296772 94654
rect 296720 94590 296772 94596
rect 295984 4004 296036 4010
rect 295984 3946 296036 3952
rect 296732 3482 296760 94590
rect 342260 94580 342312 94586
rect 342260 94522 342312 94528
rect 335358 93528 335414 93537
rect 329840 93492 329892 93498
rect 335358 93463 335414 93472
rect 329840 93434 329892 93440
rect 307760 90500 307812 90506
rect 307760 90442 307812 90448
rect 304998 84824 305054 84833
rect 304998 84759 305054 84768
rect 302240 41064 302292 41070
rect 302240 41006 302292 41012
rect 299480 28348 299532 28354
rect 299480 28290 299532 28296
rect 299492 16574 299520 28290
rect 299492 16546 300256 16574
rect 296812 10532 296864 10538
rect 296812 10474 296864 10480
rect 296824 4078 296852 10474
rect 299112 5228 299164 5234
rect 299112 5170 299164 5176
rect 296812 4072 296864 4078
rect 296812 4014 296864 4020
rect 298008 4072 298060 4078
rect 298008 4014 298060 4020
rect 296732 3454 296944 3482
rect 296916 480 296944 3454
rect 298020 480 298048 4014
rect 299124 480 299152 5170
rect 300228 480 300256 16546
rect 301320 10464 301372 10470
rect 301320 10406 301372 10412
rect 301332 480 301360 10406
rect 302252 3398 302280 41006
rect 302332 40996 302384 41002
rect 302332 40938 302384 40944
rect 302344 16574 302372 40938
rect 305012 16574 305040 84759
rect 306378 29608 306434 29617
rect 306378 29543 306434 29552
rect 306392 16574 306420 29543
rect 302344 16546 302464 16574
rect 305012 16546 305776 16574
rect 306392 16546 306880 16574
rect 302240 3392 302292 3398
rect 302240 3334 302292 3340
rect 302436 480 302464 16546
rect 304632 10396 304684 10402
rect 304632 10338 304684 10344
rect 303528 3392 303580 3398
rect 303528 3334 303580 3340
rect 303540 480 303568 3334
rect 304644 480 304672 10338
rect 305748 480 305776 16546
rect 306852 480 306880 16546
rect 307772 3482 307800 90442
rect 310520 90432 310572 90438
rect 310520 90374 310572 90380
rect 307852 30116 307904 30122
rect 307852 30058 307904 30064
rect 307864 4078 307892 30058
rect 309140 30048 309192 30054
rect 309140 29990 309192 29996
rect 309152 16574 309180 29990
rect 310532 16574 310560 90374
rect 324320 85128 324372 85134
rect 324320 85070 324372 85076
rect 313280 82272 313332 82278
rect 313280 82214 313332 82220
rect 311900 29980 311952 29986
rect 311900 29922 311952 29928
rect 311912 16574 311940 29922
rect 309152 16546 310192 16574
rect 310532 16546 311296 16574
rect 311912 16546 312400 16574
rect 307852 4072 307904 4078
rect 307852 4014 307904 4020
rect 309048 4072 309100 4078
rect 309048 4014 309100 4020
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 4014
rect 310164 480 310192 16546
rect 311268 480 311296 16546
rect 312372 480 312400 16546
rect 313292 3398 313320 82214
rect 316040 31408 316092 31414
rect 316040 31350 316092 31356
rect 313372 29912 313424 29918
rect 313372 29854 313424 29860
rect 313384 16574 313412 29854
rect 314660 29844 314712 29850
rect 314660 29786 314712 29792
rect 314672 16574 314700 29786
rect 316052 16574 316080 31350
rect 318798 31104 318854 31113
rect 318798 31039 318854 31048
rect 313384 16546 313504 16574
rect 314672 16546 315712 16574
rect 316052 16546 316816 16574
rect 313280 3392 313332 3398
rect 313280 3334 313332 3340
rect 313476 480 313504 16546
rect 314568 3392 314620 3398
rect 314568 3334 314620 3340
rect 314580 480 314608 3334
rect 315684 480 315712 16546
rect 316788 480 316816 16546
rect 317880 12164 317932 12170
rect 317880 12106 317932 12112
rect 317892 480 317920 12106
rect 318812 3398 318840 31039
rect 322938 30968 322994 30977
rect 322938 30903 322994 30912
rect 322952 16574 322980 30903
rect 322952 16546 323440 16574
rect 322294 13288 322350 13297
rect 322294 13223 322350 13232
rect 318984 12096 319036 12102
rect 318984 12038 319036 12044
rect 318800 3392 318852 3398
rect 318800 3334 318852 3340
rect 318996 480 319024 12038
rect 321190 11656 321246 11665
rect 321190 11591 321246 11600
rect 320088 3392 320140 3398
rect 320088 3334 320140 3340
rect 320100 480 320128 3334
rect 321204 480 321232 11591
rect 322308 480 322336 13223
rect 323412 480 323440 16546
rect 324332 3482 324360 85070
rect 325700 31340 325752 31346
rect 325700 31282 325752 31288
rect 324412 29776 324464 29782
rect 324412 29718 324464 29724
rect 324424 4078 324452 29718
rect 325712 16574 325740 31282
rect 328460 29708 328512 29714
rect 328460 29650 328512 29656
rect 328472 16574 328500 29650
rect 325712 16546 326752 16574
rect 328472 16546 328960 16574
rect 324412 4072 324464 4078
rect 324412 4014 324464 4020
rect 325608 4072 325660 4078
rect 325608 4014 325660 4020
rect 324332 3454 324544 3482
rect 324516 480 324544 3454
rect 325620 480 325648 4014
rect 326724 480 326752 16546
rect 327816 12028 327868 12034
rect 327816 11970 327868 11976
rect 327828 480 327856 11970
rect 328932 480 328960 16546
rect 329852 3482 329880 93434
rect 332600 32836 332652 32842
rect 332600 32778 332652 32784
rect 332612 16574 332640 32778
rect 332612 16546 333376 16574
rect 332232 13456 332284 13462
rect 332232 13398 332284 13404
rect 329932 11960 329984 11966
rect 329932 11902 329984 11908
rect 329944 4078 329972 11902
rect 329932 4072 329984 4078
rect 329932 4014 329984 4020
rect 331128 4072 331180 4078
rect 331128 4014 331180 4020
rect 329852 3454 330064 3482
rect 330036 480 330064 3454
rect 331140 480 331168 4014
rect 332244 480 332272 13398
rect 333348 480 333376 16546
rect 334440 11892 334492 11898
rect 334440 11834 334492 11840
rect 334452 480 334480 11834
rect 335372 3398 335400 93463
rect 340880 39704 340932 39710
rect 340880 39646 340932 39652
rect 336738 39400 336794 39409
rect 336738 39335 336794 39344
rect 336752 16574 336780 39335
rect 339498 24304 339554 24313
rect 339498 24239 339554 24248
rect 339512 16574 339540 24239
rect 336752 16546 337792 16574
rect 339512 16546 340000 16574
rect 335544 13388 335596 13394
rect 335544 13330 335596 13336
rect 335360 3392 335412 3398
rect 335360 3334 335412 3340
rect 335556 480 335584 13330
rect 336648 3392 336700 3398
rect 336648 3334 336700 3340
rect 336660 480 336688 3334
rect 337764 480 337792 16546
rect 338854 13152 338910 13161
rect 338854 13087 338910 13096
rect 338868 480 338896 13087
rect 339972 480 340000 16546
rect 340892 3482 340920 39646
rect 340972 31272 341024 31278
rect 340972 31214 341024 31220
rect 340984 4078 341012 31214
rect 342272 16574 342300 94522
rect 398840 94512 398892 94518
rect 398840 94454 398892 94460
rect 346400 93424 346452 93430
rect 346400 93366 346452 93372
rect 356058 93392 356114 93401
rect 345020 83496 345072 83502
rect 345020 83438 345072 83444
rect 345032 16574 345060 83438
rect 342272 16546 343312 16574
rect 345032 16546 345520 16574
rect 340972 4072 341024 4078
rect 340972 4014 341024 4020
rect 342168 4072 342220 4078
rect 342168 4014 342220 4020
rect 340892 3454 341104 3482
rect 341076 480 341104 3454
rect 342180 480 342208 4014
rect 343284 480 343312 16546
rect 344376 13320 344428 13326
rect 344376 13262 344428 13268
rect 344388 480 344416 13262
rect 345492 480 345520 16546
rect 346412 3482 346440 93366
rect 349160 93356 349212 93362
rect 356058 93327 356114 93336
rect 349160 93298 349212 93304
rect 349172 16574 349200 93298
rect 354680 31204 354732 31210
rect 354680 31146 354732 31152
rect 351918 24168 351974 24177
rect 351918 24103 351974 24112
rect 349172 16546 349936 16574
rect 346492 13252 346544 13258
rect 346492 13194 346544 13200
rect 346504 4078 346532 13194
rect 348792 11824 348844 11830
rect 348792 11766 348844 11772
rect 346492 4072 346544 4078
rect 346492 4014 346544 4020
rect 347688 4072 347740 4078
rect 347688 4014 347740 4020
rect 346412 3454 346624 3482
rect 346596 480 346624 3454
rect 347700 480 347728 4014
rect 348804 480 348832 11766
rect 349908 480 349936 16546
rect 351000 13184 351052 13190
rect 351000 13126 351052 13132
rect 351012 480 351040 13126
rect 351932 3398 351960 24103
rect 354692 16574 354720 31146
rect 356072 16574 356100 93327
rect 374000 93288 374052 93294
rect 368478 93256 368534 93265
rect 374000 93230 374052 93236
rect 368478 93191 368534 93200
rect 357440 92064 357492 92070
rect 357440 92006 357492 92012
rect 354692 16546 355456 16574
rect 356072 16546 356560 16574
rect 352104 14816 352156 14822
rect 352104 14758 352156 14764
rect 351920 3392 351972 3398
rect 351920 3334 351972 3340
rect 352116 480 352144 14758
rect 354310 13016 354366 13025
rect 354310 12951 354366 12960
rect 353208 3392 353260 3398
rect 353208 3334 353260 3340
rect 353220 480 353248 3334
rect 354324 480 354352 12951
rect 355428 480 355456 16546
rect 356532 480 356560 16546
rect 357452 3482 357480 92006
rect 362960 91996 363012 92002
rect 362960 91938 363012 91944
rect 360200 88120 360252 88126
rect 360200 88062 360252 88068
rect 357532 28280 357584 28286
rect 357532 28222 357584 28228
rect 357544 4078 357572 28222
rect 358820 24200 358872 24206
rect 358820 24142 358872 24148
rect 358832 16574 358860 24142
rect 360212 16574 360240 88062
rect 361580 31136 361632 31142
rect 361580 31078 361632 31084
rect 361592 16574 361620 31078
rect 358832 16546 359872 16574
rect 360212 16546 360976 16574
rect 361592 16546 362080 16574
rect 357532 4072 357584 4078
rect 357532 4014 357584 4020
rect 358728 4072 358780 4078
rect 358728 4014 358780 4020
rect 357452 3454 357664 3482
rect 357636 480 357664 3454
rect 358740 480 358768 4014
rect 359844 480 359872 16546
rect 360948 480 360976 16546
rect 362052 480 362080 16546
rect 362972 3398 363000 91938
rect 363052 34332 363104 34338
rect 363052 34274 363104 34280
rect 363064 16574 363092 34274
rect 365720 34264 365772 34270
rect 365720 34206 365772 34212
rect 364340 31068 364392 31074
rect 364340 31010 364392 31016
rect 364352 16574 364380 31010
rect 365732 16574 365760 34206
rect 363064 16546 363184 16574
rect 364352 16546 365392 16574
rect 365732 16546 366496 16574
rect 362960 3392 363012 3398
rect 362960 3334 363012 3340
rect 363156 480 363184 16546
rect 364248 3392 364300 3398
rect 364248 3334 364300 3340
rect 364260 480 364288 3334
rect 365364 480 365392 16546
rect 366468 480 366496 16546
rect 367560 13116 367612 13122
rect 367560 13058 367612 13064
rect 367572 480 367600 13058
rect 368492 3398 368520 93191
rect 372618 36952 372674 36961
rect 372618 36887 372674 36896
rect 372632 16574 372660 36887
rect 372632 16546 373120 16574
rect 370870 14920 370926 14929
rect 370870 14855 370926 14864
rect 368664 14748 368716 14754
rect 368664 14690 368716 14696
rect 368480 3392 368532 3398
rect 368480 3334 368532 3340
rect 368676 480 368704 14690
rect 369768 3392 369820 3398
rect 369768 3334 369820 3340
rect 369780 480 369808 3334
rect 370884 480 370912 14855
rect 371974 14784 372030 14793
rect 371974 14719 372030 14728
rect 371988 480 372016 14719
rect 373092 480 373120 16546
rect 374012 3398 374040 93230
rect 391940 93220 391992 93226
rect 391940 93162 391992 93168
rect 389178 93120 389234 93129
rect 389178 93055 389234 93064
rect 376760 85060 376812 85066
rect 376760 85002 376812 85008
rect 374092 39636 374144 39642
rect 374092 39578 374144 39584
rect 374104 16574 374132 39578
rect 375380 25764 375432 25770
rect 375380 25706 375432 25712
rect 375392 16574 375420 25706
rect 376772 16574 376800 85002
rect 379520 84992 379572 84998
rect 379520 84934 379572 84940
rect 378140 32768 378192 32774
rect 378140 32710 378192 32716
rect 378152 16574 378180 32710
rect 374104 16546 374224 16574
rect 375392 16546 376432 16574
rect 376772 16546 377536 16574
rect 378152 16546 378640 16574
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374196 480 374224 16546
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 376404 480 376432 16546
rect 377508 480 377536 16546
rect 378612 480 378640 16546
rect 379532 3398 379560 84934
rect 385038 36816 385094 36825
rect 385038 36751 385094 36760
rect 380900 32700 380952 32706
rect 380900 32642 380952 32648
rect 379612 25696 379664 25702
rect 379612 25638 379664 25644
rect 379624 16574 379652 25638
rect 380912 16574 380940 32642
rect 382280 25628 382332 25634
rect 382280 25570 382332 25576
rect 382292 16574 382320 25570
rect 379624 16546 379744 16574
rect 380912 16546 381952 16574
rect 382292 16546 383056 16574
rect 379520 3392 379572 3398
rect 379520 3334 379572 3340
rect 379716 480 379744 16546
rect 380808 3392 380860 3398
rect 380808 3334 380860 3340
rect 380820 480 380848 3334
rect 381924 480 381952 16546
rect 383028 480 383056 16546
rect 384120 14680 384172 14686
rect 384120 14622 384172 14628
rect 384132 480 384160 14622
rect 385052 3398 385080 36751
rect 385132 32632 385184 32638
rect 385132 32574 385184 32580
rect 385144 16574 385172 32574
rect 389192 16574 389220 93055
rect 390560 82204 390612 82210
rect 390560 82146 390612 82152
rect 385144 16546 385264 16574
rect 389192 16546 389680 16574
rect 385040 3392 385092 3398
rect 385040 3334 385092 3340
rect 385236 480 385264 16546
rect 387430 14648 387486 14657
rect 387430 14583 387486 14592
rect 386328 3392 386380 3398
rect 386328 3334 386380 3340
rect 386340 480 386368 3334
rect 387444 480 387472 14583
rect 388534 14512 388590 14521
rect 388534 14447 388590 14456
rect 388548 480 388576 14447
rect 389652 480 389680 16546
rect 390572 3482 390600 82146
rect 390652 32564 390704 32570
rect 390652 32506 390704 32512
rect 390664 4078 390692 32506
rect 391952 16574 391980 93162
rect 394700 32496 394752 32502
rect 394700 32438 394752 32444
rect 394712 16574 394740 32438
rect 397460 32428 397512 32434
rect 397460 32370 397512 32376
rect 396080 25560 396132 25566
rect 396080 25502 396132 25508
rect 391952 16546 392992 16574
rect 394712 16546 395200 16574
rect 390652 4072 390704 4078
rect 390652 4014 390704 4020
rect 391848 4072 391900 4078
rect 391848 4014 391900 4020
rect 390572 3454 390784 3482
rect 390756 480 390784 3454
rect 391860 480 391888 4014
rect 392964 480 392992 16546
rect 394056 14612 394108 14618
rect 394056 14554 394108 14560
rect 394068 480 394096 14554
rect 395172 480 395200 16546
rect 396092 3482 396120 25502
rect 397472 16574 397500 32370
rect 398852 16574 398880 94454
rect 401600 93152 401652 93158
rect 401600 93094 401652 93100
rect 397472 16546 398512 16574
rect 398852 16546 399616 16574
rect 396172 14544 396224 14550
rect 396172 14486 396224 14492
rect 396184 4078 396212 14486
rect 396172 4072 396224 4078
rect 396172 4014 396224 4020
rect 397368 4072 397420 4078
rect 397368 4014 397420 4020
rect 396092 3454 396304 3482
rect 396276 480 396304 3454
rect 397380 480 397408 4014
rect 398484 480 398512 16546
rect 399588 480 399616 16546
rect 400680 14476 400732 14482
rect 400680 14418 400732 14424
rect 400692 480 400720 14418
rect 401612 3398 401640 93094
rect 445760 91928 445812 91934
rect 445760 91870 445812 91876
rect 420918 90808 420974 90817
rect 420918 90743 420974 90752
rect 409880 89072 409932 89078
rect 409880 89014 409932 89020
rect 407120 87984 407172 87990
rect 407120 87926 407172 87932
rect 405738 33824 405794 33833
rect 405738 33759 405794 33768
rect 401690 32600 401746 32609
rect 401690 32535 401746 32544
rect 401704 16574 401732 32535
rect 405752 16574 405780 33759
rect 401704 16546 401824 16574
rect 405752 16546 406240 16574
rect 401600 3392 401652 3398
rect 401600 3334 401652 3340
rect 401796 480 401824 16546
rect 403990 16144 404046 16153
rect 403990 16079 404046 16088
rect 402888 3392 402940 3398
rect 402888 3334 402940 3340
rect 402900 480 402928 3334
rect 404004 480 404032 16079
rect 405094 16008 405150 16017
rect 405094 15943 405150 15952
rect 405108 480 405136 15943
rect 406212 480 406240 16546
rect 407132 3482 407160 87926
rect 408500 36576 408552 36582
rect 408500 36518 408552 36524
rect 407212 34196 407264 34202
rect 407212 34138 407264 34144
rect 407224 4078 407252 34138
rect 408512 16574 408540 36518
rect 409892 16574 409920 89014
rect 415400 38140 415452 38146
rect 415400 38082 415452 38088
rect 411260 34128 411312 34134
rect 411260 34070 411312 34076
rect 411272 16574 411300 34070
rect 414020 34060 414072 34066
rect 414020 34002 414072 34008
rect 414032 16574 414060 34002
rect 415412 16574 415440 38082
rect 418160 35488 418212 35494
rect 418160 35430 418212 35436
rect 408512 16546 409552 16574
rect 409892 16546 410656 16574
rect 411272 16546 411760 16574
rect 414032 16546 415072 16574
rect 415412 16546 416176 16574
rect 407212 4072 407264 4078
rect 407212 4014 407264 4020
rect 408408 4072 408460 4078
rect 408408 4014 408460 4020
rect 407132 3454 407344 3482
rect 407316 480 407344 3454
rect 408420 480 408448 4014
rect 409524 480 409552 16546
rect 410628 480 410656 16546
rect 411732 480 411760 16546
rect 412732 16244 412784 16250
rect 412732 16186 412784 16192
rect 412744 3398 412772 16186
rect 412824 3868 412876 3874
rect 412824 3810 412876 3816
rect 412732 3392 412784 3398
rect 412732 3334 412784 3340
rect 412836 480 412864 3810
rect 413928 3392 413980 3398
rect 413928 3334 413980 3340
rect 413940 480 413968 3334
rect 415044 480 415072 16546
rect 416148 480 416176 16546
rect 417240 16176 417292 16182
rect 417240 16118 417292 16124
rect 417252 480 417280 16118
rect 418172 3398 418200 35430
rect 420932 16574 420960 90743
rect 436098 90672 436154 90681
rect 436098 90607 436154 90616
rect 429200 89004 429252 89010
rect 429200 88946 429252 88952
rect 426440 84924 426492 84930
rect 426440 84866 426492 84872
rect 423680 40928 423732 40934
rect 423680 40870 423732 40876
rect 422300 38072 422352 38078
rect 422300 38014 422352 38020
rect 422312 16574 422340 38014
rect 420932 16546 421696 16574
rect 422312 16546 422800 16574
rect 418344 16108 418396 16114
rect 418344 16050 418396 16056
rect 418160 3392 418212 3398
rect 418160 3334 418212 3340
rect 418356 480 418384 16050
rect 420550 15872 420606 15881
rect 420550 15807 420606 15816
rect 419448 3392 419500 3398
rect 419448 3334 419500 3340
rect 419460 480 419488 3334
rect 420564 480 420592 15807
rect 421668 480 421696 16546
rect 422772 480 422800 16546
rect 423692 3482 423720 40870
rect 425060 38004 425112 38010
rect 425060 37946 425112 37952
rect 425072 16574 425100 37946
rect 426452 16574 426480 84866
rect 427820 33992 427872 33998
rect 427820 33934 427872 33940
rect 427832 16574 427860 33934
rect 425072 16546 426112 16574
rect 426452 16546 427216 16574
rect 427832 16546 428320 16574
rect 423772 16040 423824 16046
rect 423772 15982 423824 15988
rect 423784 3874 423812 15982
rect 423772 3868 423824 3874
rect 423772 3810 423824 3816
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 423692 3454 423904 3482
rect 423876 480 423904 3454
rect 424980 480 425008 3810
rect 426084 480 426112 16546
rect 427188 480 427216 16546
rect 428292 480 428320 16546
rect 429212 3398 429240 88946
rect 429292 87916 429344 87922
rect 429292 87858 429344 87864
rect 429304 16574 429332 87858
rect 433340 86352 433392 86358
rect 433340 86294 433392 86300
rect 431960 37936 432012 37942
rect 431960 37878 432012 37884
rect 430580 33924 430632 33930
rect 430580 33866 430632 33872
rect 430592 16574 430620 33866
rect 431972 16574 432000 37878
rect 433352 16574 433380 86294
rect 434720 80776 434772 80782
rect 434720 80718 434772 80724
rect 429304 16546 429424 16574
rect 430592 16546 431632 16574
rect 431972 16546 432736 16574
rect 433352 16546 433840 16574
rect 429200 3392 429252 3398
rect 429200 3334 429252 3340
rect 429396 480 429424 16546
rect 430488 3392 430540 3398
rect 430488 3334 430540 3340
rect 430500 480 430528 3334
rect 431604 480 431632 16546
rect 432708 480 432736 16546
rect 433812 480 433840 16546
rect 434732 3398 434760 80718
rect 434810 35728 434866 35737
rect 434810 35663 434866 35672
rect 434824 16574 434852 35663
rect 436112 16574 436140 90607
rect 440240 84856 440292 84862
rect 440240 84798 440292 84804
rect 438858 38040 438914 38049
rect 438858 37975 438914 37984
rect 437478 35592 437534 35601
rect 437478 35527 437534 35536
rect 437492 16574 437520 35527
rect 438872 16574 438900 37975
rect 434824 16546 434944 16574
rect 436112 16546 437152 16574
rect 437492 16546 438256 16574
rect 438872 16546 439360 16574
rect 434720 3392 434772 3398
rect 434720 3334 434772 3340
rect 434916 480 434944 16546
rect 436008 3392 436060 3398
rect 436008 3334 436060 3340
rect 436020 480 436048 3334
rect 437124 480 437152 16546
rect 438228 480 438256 16546
rect 439332 480 439360 16546
rect 440252 3482 440280 84798
rect 443000 39568 443052 39574
rect 443000 39510 443052 39516
rect 440332 35420 440384 35426
rect 440332 35362 440384 35368
rect 440344 3874 440372 35362
rect 443012 16574 443040 39510
rect 444380 35352 444432 35358
rect 444380 35294 444432 35300
rect 444392 16574 444420 35294
rect 443012 16546 443776 16574
rect 444392 16546 444880 16574
rect 440332 3868 440384 3874
rect 440332 3810 440384 3816
rect 441528 3868 441580 3874
rect 441528 3810 441580 3816
rect 440252 3454 440464 3482
rect 440436 480 440464 3454
rect 441540 480 441568 3810
rect 442632 3800 442684 3806
rect 442632 3742 442684 3748
rect 442644 480 442672 3742
rect 443748 480 443776 16546
rect 444852 480 444880 16546
rect 445772 3482 445800 91870
rect 445852 86284 445904 86290
rect 445852 86226 445904 86232
rect 445864 3806 445892 86226
rect 446416 3874 446444 97242
rect 498200 96144 498252 96150
rect 471978 96112 472034 96121
rect 498200 96086 498252 96092
rect 471978 96047 472034 96056
rect 456800 91860 456852 91866
rect 456800 91802 456852 91808
rect 448520 53168 448572 53174
rect 448520 53110 448572 53116
rect 447140 33856 447192 33862
rect 447140 33798 447192 33804
rect 447152 16574 447180 33798
rect 448532 16574 448560 53110
rect 455420 53100 455472 53106
rect 455420 53042 455472 53048
rect 451278 37904 451334 37913
rect 451278 37839 451334 37848
rect 449898 17504 449954 17513
rect 449898 17439 449954 17448
rect 449912 16574 449940 17439
rect 447152 16546 448192 16574
rect 448532 16546 449296 16574
rect 449912 16546 450400 16574
rect 446404 3868 446456 3874
rect 446404 3810 446456 3816
rect 445852 3800 445904 3806
rect 445852 3742 445904 3748
rect 447048 3800 447100 3806
rect 447048 3742 447100 3748
rect 445772 3454 445984 3482
rect 445956 480 445984 3454
rect 447060 480 447088 3742
rect 448164 480 448192 16546
rect 449268 480 449296 16546
rect 450372 480 450400 16546
rect 451292 3398 451320 37839
rect 451370 35456 451426 35465
rect 451370 35391 451426 35400
rect 451384 16574 451412 35391
rect 454038 35320 454094 35329
rect 454038 35255 454094 35264
rect 452658 17368 452714 17377
rect 452658 17303 452714 17312
rect 452672 16574 452700 17303
rect 454052 16574 454080 35255
rect 455432 16574 455460 53042
rect 451384 16546 451504 16574
rect 452672 16546 453712 16574
rect 454052 16546 454816 16574
rect 455432 16546 455920 16574
rect 451280 3392 451332 3398
rect 451280 3334 451332 3340
rect 451476 480 451504 16546
rect 452568 3392 452620 3398
rect 452568 3334 452620 3340
rect 452580 480 452608 3334
rect 453684 480 453712 16546
rect 454788 480 454816 16546
rect 455892 480 455920 16546
rect 456708 3732 456760 3738
rect 456708 3674 456760 3680
rect 456720 3398 456748 3674
rect 456812 3482 456840 91802
rect 469220 88052 469272 88058
rect 469220 87994 469272 88000
rect 462320 54528 462372 54534
rect 462320 54470 462372 54476
rect 456892 40860 456944 40866
rect 456892 40802 456944 40808
rect 456904 3738 456932 40802
rect 460940 40792 460992 40798
rect 460940 40734 460992 40740
rect 459560 17536 459612 17542
rect 459560 17478 459612 17484
rect 459572 16574 459600 17478
rect 460952 16574 460980 40734
rect 459572 16546 460336 16574
rect 460952 16546 461440 16574
rect 456892 3732 456944 3738
rect 456892 3674 456944 3680
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 456812 3454 457024 3482
rect 456708 3392 456760 3398
rect 456708 3334 456760 3340
rect 456996 480 457024 3454
rect 458100 480 458128 3674
rect 459192 3392 459244 3398
rect 459192 3334 459244 3340
rect 459204 480 459232 3334
rect 460308 480 460336 16546
rect 461412 480 461440 16546
rect 462332 3482 462360 54470
rect 465080 40724 465132 40730
rect 465080 40666 465132 40672
rect 463700 24132 463752 24138
rect 463700 24074 463752 24080
rect 462412 17468 462464 17474
rect 462412 17410 462464 17416
rect 462424 3738 462452 17410
rect 463712 16574 463740 24074
rect 465092 16574 465120 40666
rect 467930 32464 467986 32473
rect 467930 32399 467986 32408
rect 466460 18828 466512 18834
rect 466460 18770 466512 18776
rect 466472 16574 466500 18770
rect 467944 16574 467972 32399
rect 469232 16574 469260 87994
rect 470598 18864 470654 18873
rect 470598 18799 470654 18808
rect 470612 16574 470640 18799
rect 471992 16574 472020 96047
rect 488538 95976 488594 95985
rect 488538 95911 488594 95920
rect 485778 90536 485834 90545
rect 485778 90471 485834 90480
rect 473452 90364 473504 90370
rect 473452 90306 473504 90312
rect 463712 16546 464752 16574
rect 465092 16546 465856 16574
rect 466472 16546 466960 16574
rect 467944 16546 468064 16574
rect 469232 16546 470272 16574
rect 470612 16546 471376 16574
rect 471992 16546 472480 16574
rect 462412 3732 462464 3738
rect 462412 3674 462464 3680
rect 463608 3732 463660 3738
rect 463608 3674 463660 3680
rect 462332 3454 462544 3482
rect 462516 480 462544 3454
rect 463620 480 463648 3674
rect 464724 480 464752 16546
rect 465828 480 465856 16546
rect 466932 480 466960 16546
rect 468036 480 468064 16546
rect 469128 4004 469180 4010
rect 469128 3946 469180 3952
rect 469140 480 469168 3946
rect 470244 480 470272 16546
rect 471348 480 471376 16546
rect 472452 480 472480 16546
rect 473464 3602 473492 90306
rect 483020 39500 483072 39506
rect 483020 39442 483072 39448
rect 478880 35284 478932 35290
rect 478880 35226 478932 35232
rect 477500 18760 477552 18766
rect 477500 18702 477552 18708
rect 474740 17400 474792 17406
rect 474740 17342 474792 17348
rect 474752 16574 474780 17342
rect 477512 16574 477540 18702
rect 474752 16546 475792 16574
rect 477512 16546 478000 16574
rect 473544 3664 473596 3670
rect 473544 3606 473596 3612
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 473556 480 473584 3606
rect 474648 3596 474700 3602
rect 474648 3538 474700 3544
rect 474660 480 474688 3538
rect 475764 480 475792 16546
rect 476856 3732 476908 3738
rect 476856 3674 476908 3680
rect 476868 480 476896 3674
rect 477972 480 478000 16546
rect 478892 1154 478920 35226
rect 481640 33788 481692 33794
rect 481640 33730 481692 33736
rect 478972 29640 479024 29646
rect 478972 29582 479024 29588
rect 478984 16574 479012 29582
rect 481652 16574 481680 33730
rect 483032 16574 483060 39442
rect 484398 35184 484454 35193
rect 484398 35119 484454 35128
rect 478984 16546 479104 16574
rect 481652 16546 482416 16574
rect 483032 16546 483520 16574
rect 478880 1148 478932 1154
rect 478880 1090 478932 1096
rect 479076 480 479104 16546
rect 481272 5160 481324 5166
rect 481272 5102 481324 5108
rect 480168 1148 480220 1154
rect 480168 1090 480220 1096
rect 480180 480 480208 1090
rect 481284 480 481312 5102
rect 482388 480 482416 16546
rect 483492 480 483520 16546
rect 484412 3602 484440 35119
rect 485792 16574 485820 90471
rect 488552 16574 488580 95911
rect 490012 20392 490064 20398
rect 490012 20334 490064 20340
rect 485792 16546 486832 16574
rect 488552 16546 489040 16574
rect 484582 6488 484638 6497
rect 484582 6423 484638 6432
rect 484400 3596 484452 3602
rect 484400 3538 484452 3544
rect 484596 480 484624 6423
rect 485688 3596 485740 3602
rect 485688 3538 485740 3544
rect 485700 480 485728 3538
rect 486804 480 486832 16546
rect 487894 6352 487950 6361
rect 487894 6287 487950 6296
rect 487908 480 487936 6287
rect 489012 480 489040 16546
rect 490024 3534 490052 20334
rect 494060 20324 494112 20330
rect 494060 20266 494112 20272
rect 491300 17332 491352 17338
rect 491300 17274 491352 17280
rect 491312 16574 491340 17274
rect 494072 16574 494100 20266
rect 496820 20256 496872 20262
rect 496820 20198 496872 20204
rect 495532 17264 495584 17270
rect 495532 17206 495584 17212
rect 495544 16574 495572 17206
rect 496832 16574 496860 20198
rect 498212 16574 498240 96086
rect 514760 96076 514812 96082
rect 514760 96018 514812 96024
rect 506480 91792 506532 91798
rect 506480 91734 506532 91740
rect 502338 90400 502394 90409
rect 502338 90335 502394 90344
rect 500960 20188 501012 20194
rect 500960 20130 501012 20136
rect 491312 16546 492352 16574
rect 494072 16546 494560 16574
rect 495544 16546 495664 16574
rect 496832 16546 497872 16574
rect 498212 16546 498976 16574
rect 490104 3936 490156 3942
rect 490104 3878 490156 3884
rect 490012 3528 490064 3534
rect 490012 3470 490064 3476
rect 490116 480 490144 3878
rect 491208 3528 491260 3534
rect 491208 3470 491260 3476
rect 491220 480 491248 3470
rect 492324 480 492352 16546
rect 493416 3596 493468 3602
rect 493416 3538 493468 3544
rect 493428 480 493456 3538
rect 494532 480 494560 16546
rect 495636 480 495664 16546
rect 496728 3460 496780 3466
rect 496728 3402 496780 3408
rect 496740 480 496768 3402
rect 497844 480 497872 16546
rect 498948 480 498976 16546
rect 500040 5092 500092 5098
rect 500040 5034 500092 5040
rect 500052 480 500080 5034
rect 500972 3482 501000 20130
rect 501050 17232 501106 17241
rect 501050 17167 501106 17176
rect 501064 3602 501092 17167
rect 502352 16574 502380 90335
rect 505098 18728 505154 18737
rect 505098 18663 505154 18672
rect 505112 16574 505140 18663
rect 502352 16546 503392 16574
rect 505112 16546 505600 16574
rect 501052 3596 501104 3602
rect 501052 3538 501104 3544
rect 502248 3596 502300 3602
rect 502248 3538 502300 3544
rect 500972 3454 501184 3482
rect 501156 480 501184 3454
rect 502260 480 502288 3538
rect 503364 480 503392 16546
rect 504454 6216 504510 6225
rect 504454 6151 504510 6160
rect 504468 480 504496 6151
rect 505572 480 505600 16546
rect 506492 3482 506520 91734
rect 512000 87848 512052 87854
rect 512000 87790 512052 87796
rect 507860 80708 507912 80714
rect 507860 80650 507912 80656
rect 506572 21684 506624 21690
rect 506572 21626 506624 21632
rect 506584 3602 506612 21626
rect 507872 16574 507900 80650
rect 510620 21616 510672 21622
rect 510620 21558 510672 21564
rect 510632 16574 510660 21558
rect 507872 16546 508912 16574
rect 510632 16546 511120 16574
rect 506572 3596 506624 3602
rect 506572 3538 506624 3544
rect 507768 3596 507820 3602
rect 507768 3538 507820 3544
rect 506492 3454 506704 3482
rect 506676 480 506704 3454
rect 507780 480 507808 3538
rect 508884 480 508912 16546
rect 509976 5024 510028 5030
rect 509976 4966 510028 4972
rect 509988 480 510016 4966
rect 511092 480 511120 16546
rect 512012 3534 512040 87790
rect 512092 82136 512144 82142
rect 512092 82078 512144 82084
rect 512104 16574 512132 82078
rect 513380 21548 513432 21554
rect 513380 21490 513432 21496
rect 513392 16574 513420 21490
rect 514772 16574 514800 96018
rect 528560 96008 528612 96014
rect 528560 95950 528612 95956
rect 521658 95840 521714 95849
rect 521658 95775 521714 95784
rect 516140 87780 516192 87786
rect 516140 87722 516192 87728
rect 516152 16574 516180 87722
rect 520278 21312 520334 21321
rect 520278 21247 520334 21256
rect 517520 18692 517572 18698
rect 517520 18634 517572 18640
rect 512104 16546 512224 16574
rect 513392 16546 514432 16574
rect 514772 16546 515536 16574
rect 516152 16546 516640 16574
rect 512000 3528 512052 3534
rect 512000 3470 512052 3476
rect 512196 480 512224 16546
rect 513288 3528 513340 3534
rect 513288 3470 513340 3476
rect 513300 480 513328 3470
rect 514404 480 514432 16546
rect 515508 480 515536 16546
rect 516612 480 516640 16546
rect 517532 7546 517560 18634
rect 520292 16574 520320 21247
rect 521672 16574 521700 95775
rect 523132 21480 523184 21486
rect 523132 21422 523184 21428
rect 520292 16546 521056 16574
rect 521672 16546 522160 16574
rect 517520 7540 517572 7546
rect 517520 7482 517572 7488
rect 518808 7540 518860 7546
rect 518808 7482 518860 7488
rect 517704 6384 517756 6390
rect 517704 6326 517756 6332
rect 516784 4888 516836 4894
rect 516784 4830 516836 4836
rect 516796 4758 516824 4830
rect 516784 4752 516836 4758
rect 516784 4694 516836 4700
rect 517716 480 517744 6326
rect 518820 480 518848 7482
rect 519910 4856 519966 4865
rect 519910 4791 519966 4800
rect 519924 480 519952 4791
rect 521028 480 521056 16546
rect 522132 480 522160 16546
rect 523144 7546 523172 21422
rect 524420 18624 524472 18630
rect 524420 18566 524472 18572
rect 524432 16574 524460 18566
rect 528572 16574 528600 95950
rect 545120 95940 545172 95946
rect 545120 95882 545172 95888
rect 535458 79384 535514 79393
rect 535458 79319 535514 79328
rect 532700 39432 532752 39438
rect 532700 39374 532752 39380
rect 531320 35216 531372 35222
rect 531320 35158 531372 35164
rect 531332 16574 531360 35158
rect 532712 16574 532740 39374
rect 534078 18592 534134 18601
rect 534078 18527 534134 18536
rect 524432 16546 525472 16574
rect 528572 16546 528784 16574
rect 531332 16546 532096 16574
rect 532712 16546 533200 16574
rect 523132 7540 523184 7546
rect 523132 7482 523184 7488
rect 524328 7540 524380 7546
rect 524328 7482 524380 7488
rect 523224 3800 523276 3806
rect 523224 3742 523276 3748
rect 523236 480 523264 3742
rect 524340 480 524368 7482
rect 525444 480 525472 16546
rect 527640 7744 527692 7750
rect 527640 7686 527692 7692
rect 526536 4956 526588 4962
rect 526536 4898 526588 4904
rect 526548 480 526576 4898
rect 527652 480 527680 7686
rect 528756 480 528784 16546
rect 530952 7676 531004 7682
rect 530952 7618 531004 7624
rect 529848 4752 529900 4758
rect 529848 4694 529900 4700
rect 529860 480 529888 4694
rect 530964 480 530992 7618
rect 532068 480 532096 16546
rect 533172 480 533200 16546
rect 534092 746 534120 18527
rect 535472 16574 535500 79319
rect 542360 39364 542412 39370
rect 542360 39306 542412 39312
rect 538218 36680 538274 36689
rect 538218 36615 538274 36624
rect 536838 22808 536894 22817
rect 536838 22743 536894 22752
rect 536852 16574 536880 22743
rect 538232 16574 538260 36615
rect 542372 16574 542400 39306
rect 535472 16546 536512 16574
rect 536852 16546 537616 16574
rect 538232 16546 538720 16574
rect 542372 16546 543136 16574
rect 534264 7608 534316 7614
rect 534264 7550 534316 7556
rect 534080 740 534132 746
rect 534080 682 534132 688
rect 534276 480 534304 7550
rect 535368 740 535420 746
rect 535368 682 535420 688
rect 535380 480 535408 682
rect 536484 480 536512 16546
rect 537588 480 537616 16546
rect 538692 480 538720 16546
rect 541992 15972 542044 15978
rect 541992 15914 542044 15920
rect 539600 10328 539652 10334
rect 539600 10270 539652 10276
rect 539612 3534 539640 10270
rect 539784 6316 539836 6322
rect 539784 6258 539836 6264
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539796 480 539824 6258
rect 540888 3528 540940 3534
rect 540888 3470 540940 3476
rect 540900 480 540928 3470
rect 542004 480 542032 15914
rect 543108 480 543136 16546
rect 544200 11756 544252 11762
rect 544200 11698 544252 11704
rect 544212 480 544240 11698
rect 545132 3482 545160 95882
rect 545212 87712 545264 87718
rect 545212 87654 545264 87660
rect 545224 3602 545252 87654
rect 549260 87644 549312 87650
rect 549260 87586 549312 87592
rect 546500 20120 546552 20126
rect 546500 20062 546552 20068
rect 546512 16574 546540 20062
rect 549272 16574 549300 87586
rect 579620 71732 579672 71738
rect 579620 71674 579672 71680
rect 579632 70417 579660 71674
rect 579618 70408 579674 70417
rect 579618 70343 579674 70352
rect 552018 39264 552074 39273
rect 552018 39199 552074 39208
rect 550640 21412 550692 21418
rect 550640 21354 550692 21360
rect 546512 16546 547552 16574
rect 549272 16546 549760 16574
rect 545212 3596 545264 3602
rect 545212 3538 545264 3544
rect 546408 3596 546460 3602
rect 546408 3538 546460 3544
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546420 480 546448 3538
rect 547524 480 547552 16546
rect 548616 4820 548668 4826
rect 548616 4762 548668 4768
rect 548628 480 548656 4762
rect 549732 480 549760 16546
rect 550652 3482 550680 21354
rect 550730 19952 550786 19961
rect 550730 19887 550786 19896
rect 550744 3602 550772 19887
rect 552032 16574 552060 39199
rect 554778 36544 554834 36553
rect 554778 36479 554834 36488
rect 553398 22672 553454 22681
rect 553398 22607 553454 22616
rect 553412 16574 553440 22607
rect 554792 16574 554820 36479
rect 557540 20052 557592 20058
rect 557540 19994 557592 20000
rect 557552 16574 557580 19994
rect 561680 19984 561732 19990
rect 561680 19926 561732 19932
rect 561692 16574 561720 19926
rect 552032 16546 553072 16574
rect 553412 16546 554176 16574
rect 554792 16546 555280 16574
rect 557552 16546 558592 16574
rect 561692 16546 561904 16574
rect 550732 3596 550784 3602
rect 550732 3538 550784 3544
rect 551928 3596 551980 3602
rect 551928 3538 551980 3544
rect 550652 3454 550864 3482
rect 550836 480 550864 3454
rect 551940 480 551968 3538
rect 553044 480 553072 16546
rect 554148 480 554176 16546
rect 555252 480 555280 16546
rect 557448 8968 557500 8974
rect 557448 8910 557500 8916
rect 556344 6248 556396 6254
rect 556344 6190 556396 6196
rect 556356 480 556384 6190
rect 557460 480 557488 8910
rect 558564 480 558592 16546
rect 560760 15904 560812 15910
rect 560760 15846 560812 15852
rect 559656 6180 559708 6186
rect 559656 6122 559708 6128
rect 559668 480 559696 6122
rect 560772 480 560800 15846
rect 561876 480 561904 16546
rect 580276 7857 580304 149398
rect 580368 23497 580396 151030
rect 580632 149320 580684 149326
rect 580632 149262 580684 149268
rect 580540 149252 580592 149258
rect 580540 149194 580592 149200
rect 580448 149184 580500 149190
rect 580448 149126 580500 149132
rect 580460 54777 580488 149126
rect 580552 86057 580580 149194
rect 580644 101697 580672 149262
rect 580630 101688 580686 101697
rect 580630 101623 580686 101632
rect 580538 86048 580594 86057
rect 580538 85983 580594 85992
rect 580446 54768 580502 54777
rect 580446 54703 580502 54712
rect 580354 23488 580410 23497
rect 580354 23423 580410 23432
rect 580262 7848 580318 7857
rect 580262 7783 580318 7792
rect 87616 354 87644 462
rect 87114 326 87644 354
rect 87114 -960 87226 326
rect 88218 -960 88330 480
rect 89322 -960 89434 480
rect 90426 -960 90538 480
rect 91530 -960 91642 480
rect 92634 -960 92746 480
rect 93738 -960 93850 480
rect 94842 -960 94954 480
rect 95946 -960 96058 480
rect 97050 -960 97162 480
rect 98154 -960 98266 480
rect 99258 -960 99370 480
rect 100362 -960 100474 480
rect 101466 -960 101578 480
rect 102570 -960 102682 480
rect 103674 -960 103786 480
rect 104778 -960 104890 480
rect 105882 -960 105994 480
rect 106986 -960 107098 480
rect 108090 -960 108202 480
rect 109194 -960 109306 480
rect 110298 -960 110410 480
rect 111402 -960 111514 480
rect 112506 -960 112618 480
rect 113610 -960 113722 480
rect 114714 -960 114826 480
rect 115818 -960 115930 480
rect 116922 -960 117034 480
rect 118026 -960 118138 480
rect 119130 -960 119242 480
rect 120234 -960 120346 480
rect 121338 -960 121450 480
rect 122442 -960 122554 480
rect 123546 -960 123658 480
rect 124650 -960 124762 480
rect 125754 -960 125866 480
rect 126858 -960 126970 480
rect 127962 -960 128074 480
rect 129066 -960 129178 480
rect 130170 -960 130282 480
rect 131274 -960 131386 480
rect 132378 -960 132490 480
rect 133482 -960 133594 480
rect 134586 -960 134698 480
rect 135690 -960 135802 480
rect 136794 -960 136906 480
rect 137898 -960 138010 480
rect 139002 -960 139114 480
rect 140106 -960 140218 480
rect 141210 -960 141322 480
rect 142314 -960 142426 480
rect 143418 -960 143530 480
rect 144522 -960 144634 480
rect 145626 -960 145738 480
rect 146730 -960 146842 480
rect 147834 -960 147946 480
rect 148938 -960 149050 480
rect 150042 -960 150154 480
rect 151146 -960 151258 480
rect 152250 -960 152362 480
rect 153354 -960 153466 480
rect 154458 -960 154570 480
rect 155562 -960 155674 480
rect 156666 -960 156778 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 159978 -960 160090 480
rect 161082 -960 161194 480
rect 162186 -960 162298 480
rect 163290 -960 163402 480
rect 164394 -960 164506 480
rect 165498 -960 165610 480
rect 166602 -960 166714 480
rect 167706 -960 167818 480
rect 168810 -960 168922 480
rect 169914 -960 170026 480
rect 171018 -960 171130 480
rect 172122 -960 172234 480
rect 173226 -960 173338 480
rect 174330 -960 174442 480
rect 175434 -960 175546 480
rect 176538 -960 176650 480
rect 177642 -960 177754 480
rect 178746 -960 178858 480
rect 179850 -960 179962 480
rect 180954 -960 181066 480
rect 182058 -960 182170 480
rect 183162 -960 183274 480
rect 184266 -960 184378 480
rect 185370 -960 185482 480
rect 186474 -960 186586 480
rect 187578 -960 187690 480
rect 188682 -960 188794 480
rect 189786 -960 189898 480
rect 190890 -960 191002 480
rect 191994 -960 192106 480
rect 193098 -960 193210 480
rect 194202 -960 194314 480
rect 195306 -960 195418 480
rect 196410 -960 196522 480
rect 197514 -960 197626 480
rect 198618 -960 198730 480
rect 199722 -960 199834 480
rect 200826 -960 200938 480
rect 201930 -960 202042 480
rect 203034 -960 203146 480
rect 204138 -960 204250 480
rect 205242 -960 205354 480
rect 206346 -960 206458 480
rect 207450 -960 207562 480
rect 208554 -960 208666 480
rect 209658 -960 209770 480
rect 210762 -960 210874 480
rect 211866 -960 211978 480
rect 212970 -960 213082 480
rect 214074 -960 214186 480
rect 215178 -960 215290 480
rect 216282 -960 216394 480
rect 217386 -960 217498 480
rect 218490 -960 218602 480
rect 219594 -960 219706 480
rect 220698 -960 220810 480
rect 221802 -960 221914 480
rect 222906 -960 223018 480
rect 224010 -960 224122 480
rect 225114 -960 225226 480
rect 226218 -960 226330 480
rect 227322 -960 227434 480
rect 228426 -960 228538 480
rect 229530 -960 229642 480
rect 230634 -960 230746 480
rect 231738 -960 231850 480
rect 232842 -960 232954 480
rect 233946 -960 234058 480
rect 235050 -960 235162 480
rect 236154 -960 236266 480
rect 237258 -960 237370 480
rect 238362 -960 238474 480
rect 239466 -960 239578 480
rect 240570 -960 240682 480
rect 241674 -960 241786 480
rect 242778 -960 242890 480
rect 243882 -960 243994 480
rect 244986 -960 245098 480
rect 246090 -960 246202 480
rect 247194 -960 247306 480
rect 248298 -960 248410 480
rect 249402 -960 249514 480
rect 250506 -960 250618 480
rect 251610 -960 251722 480
rect 252714 -960 252826 480
rect 253818 -960 253930 480
rect 254922 -960 255034 480
rect 256026 -960 256138 480
rect 257130 -960 257242 480
rect 258234 -960 258346 480
rect 259338 -960 259450 480
rect 260442 -960 260554 480
rect 261546 -960 261658 480
rect 262650 -960 262762 480
rect 263754 -960 263866 480
rect 264858 -960 264970 480
rect 265962 -960 266074 480
rect 267066 -960 267178 480
rect 268170 -960 268282 480
rect 269274 -960 269386 480
rect 270378 -960 270490 480
rect 271482 -960 271594 480
rect 272586 -960 272698 480
rect 273690 -960 273802 480
rect 274794 -960 274906 480
rect 275898 -960 276010 480
rect 277002 -960 277114 480
rect 278106 -960 278218 480
rect 279210 -960 279322 480
rect 280314 -960 280426 480
rect 281418 -960 281530 480
rect 282522 -960 282634 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285834 -960 285946 480
rect 286938 -960 287050 480
rect 288042 -960 288154 480
rect 289146 -960 289258 480
rect 290250 -960 290362 480
rect 291354 -960 291466 480
rect 292458 -960 292570 480
rect 293562 -960 293674 480
rect 294666 -960 294778 480
rect 295770 -960 295882 480
rect 296874 -960 296986 480
rect 297978 -960 298090 480
rect 299082 -960 299194 480
rect 300186 -960 300298 480
rect 301290 -960 301402 480
rect 302394 -960 302506 480
rect 303498 -960 303610 480
rect 304602 -960 304714 480
rect 305706 -960 305818 480
rect 306810 -960 306922 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310122 -960 310234 480
rect 311226 -960 311338 480
rect 312330 -960 312442 480
rect 313434 -960 313546 480
rect 314538 -960 314650 480
rect 315642 -960 315754 480
rect 316746 -960 316858 480
rect 317850 -960 317962 480
rect 318954 -960 319066 480
rect 320058 -960 320170 480
rect 321162 -960 321274 480
rect 322266 -960 322378 480
rect 323370 -960 323482 480
rect 324474 -960 324586 480
rect 325578 -960 325690 480
rect 326682 -960 326794 480
rect 327786 -960 327898 480
rect 328890 -960 329002 480
rect 329994 -960 330106 480
rect 331098 -960 331210 480
rect 332202 -960 332314 480
rect 333306 -960 333418 480
rect 334410 -960 334522 480
rect 335514 -960 335626 480
rect 336618 -960 336730 480
rect 337722 -960 337834 480
rect 338826 -960 338938 480
rect 339930 -960 340042 480
rect 341034 -960 341146 480
rect 342138 -960 342250 480
rect 343242 -960 343354 480
rect 344346 -960 344458 480
rect 345450 -960 345562 480
rect 346554 -960 346666 480
rect 347658 -960 347770 480
rect 348762 -960 348874 480
rect 349866 -960 349978 480
rect 350970 -960 351082 480
rect 352074 -960 352186 480
rect 353178 -960 353290 480
rect 354282 -960 354394 480
rect 355386 -960 355498 480
rect 356490 -960 356602 480
rect 357594 -960 357706 480
rect 358698 -960 358810 480
rect 359802 -960 359914 480
rect 360906 -960 361018 480
rect 362010 -960 362122 480
rect 363114 -960 363226 480
rect 364218 -960 364330 480
rect 365322 -960 365434 480
rect 366426 -960 366538 480
rect 367530 -960 367642 480
rect 368634 -960 368746 480
rect 369738 -960 369850 480
rect 370842 -960 370954 480
rect 371946 -960 372058 480
rect 373050 -960 373162 480
rect 374154 -960 374266 480
rect 375258 -960 375370 480
rect 376362 -960 376474 480
rect 377466 -960 377578 480
rect 378570 -960 378682 480
rect 379674 -960 379786 480
rect 380778 -960 380890 480
rect 381882 -960 381994 480
rect 382986 -960 383098 480
rect 384090 -960 384202 480
rect 385194 -960 385306 480
rect 386298 -960 386410 480
rect 387402 -960 387514 480
rect 388506 -960 388618 480
rect 389610 -960 389722 480
rect 390714 -960 390826 480
rect 391818 -960 391930 480
rect 392922 -960 393034 480
rect 394026 -960 394138 480
rect 395130 -960 395242 480
rect 396234 -960 396346 480
rect 397338 -960 397450 480
rect 398442 -960 398554 480
rect 399546 -960 399658 480
rect 400650 -960 400762 480
rect 401754 -960 401866 480
rect 402858 -960 402970 480
rect 403962 -960 404074 480
rect 405066 -960 405178 480
rect 406170 -960 406282 480
rect 407274 -960 407386 480
rect 408378 -960 408490 480
rect 409482 -960 409594 480
rect 410586 -960 410698 480
rect 411690 -960 411802 480
rect 412794 -960 412906 480
rect 413898 -960 414010 480
rect 415002 -960 415114 480
rect 416106 -960 416218 480
rect 417210 -960 417322 480
rect 418314 -960 418426 480
rect 419418 -960 419530 480
rect 420522 -960 420634 480
rect 421626 -960 421738 480
rect 422730 -960 422842 480
rect 423834 -960 423946 480
rect 424938 -960 425050 480
rect 426042 -960 426154 480
rect 427146 -960 427258 480
rect 428250 -960 428362 480
rect 429354 -960 429466 480
rect 430458 -960 430570 480
rect 431562 -960 431674 480
rect 432666 -960 432778 480
rect 433770 -960 433882 480
rect 434874 -960 434986 480
rect 435978 -960 436090 480
rect 437082 -960 437194 480
rect 438186 -960 438298 480
rect 439290 -960 439402 480
rect 440394 -960 440506 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443706 -960 443818 480
rect 444810 -960 444922 480
rect 445914 -960 446026 480
rect 447018 -960 447130 480
rect 448122 -960 448234 480
rect 449226 -960 449338 480
rect 450330 -960 450442 480
rect 451434 -960 451546 480
rect 452538 -960 452650 480
rect 453642 -960 453754 480
rect 454746 -960 454858 480
rect 455850 -960 455962 480
rect 456954 -960 457066 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460266 -960 460378 480
rect 461370 -960 461482 480
rect 462474 -960 462586 480
rect 463578 -960 463690 480
rect 464682 -960 464794 480
rect 465786 -960 465898 480
rect 466890 -960 467002 480
rect 467994 -960 468106 480
rect 469098 -960 469210 480
rect 470202 -960 470314 480
rect 471306 -960 471418 480
rect 472410 -960 472522 480
rect 473514 -960 473626 480
rect 474618 -960 474730 480
rect 475722 -960 475834 480
rect 476826 -960 476938 480
rect 477930 -960 478042 480
rect 479034 -960 479146 480
rect 480138 -960 480250 480
rect 481242 -960 481354 480
rect 482346 -960 482458 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485658 -960 485770 480
rect 486762 -960 486874 480
rect 487866 -960 487978 480
rect 488970 -960 489082 480
rect 490074 -960 490186 480
rect 491178 -960 491290 480
rect 492282 -960 492394 480
rect 493386 -960 493498 480
rect 494490 -960 494602 480
rect 495594 -960 495706 480
rect 496698 -960 496810 480
rect 497802 -960 497914 480
rect 498906 -960 499018 480
rect 500010 -960 500122 480
rect 501114 -960 501226 480
rect 502218 -960 502330 480
rect 503322 -960 503434 480
rect 504426 -960 504538 480
rect 505530 -960 505642 480
rect 506634 -960 506746 480
rect 507738 -960 507850 480
rect 508842 -960 508954 480
rect 509946 -960 510058 480
rect 511050 -960 511162 480
rect 512154 -960 512266 480
rect 513258 -960 513370 480
rect 514362 -960 514474 480
rect 515466 -960 515578 480
rect 516570 -960 516682 480
rect 517674 -960 517786 480
rect 518778 -960 518890 480
rect 519882 -960 519994 480
rect 520986 -960 521098 480
rect 522090 -960 522202 480
rect 523194 -960 523306 480
rect 524298 -960 524410 480
rect 525402 -960 525514 480
rect 526506 -960 526618 480
rect 527610 -960 527722 480
rect 528714 -960 528826 480
rect 529818 -960 529930 480
rect 530922 -960 531034 480
rect 532026 -960 532138 480
rect 533130 -960 533242 480
rect 534234 -960 534346 480
rect 535338 -960 535450 480
rect 536442 -960 536554 480
rect 537546 -960 537658 480
rect 538650 -960 538762 480
rect 539754 -960 539866 480
rect 540858 -960 540970 480
rect 541962 -960 542074 480
rect 543066 -960 543178 480
rect 544170 -960 544282 480
rect 545274 -960 545386 480
rect 546378 -960 546490 480
rect 547482 -960 547594 480
rect 548586 -960 548698 480
rect 549690 -960 549802 480
rect 550794 -960 550906 480
rect 551898 -960 552010 480
rect 553002 -960 553114 480
rect 554106 -960 554218 480
rect 555210 -960 555322 480
rect 556314 -960 556426 480
rect 557418 -960 557530 480
rect 558522 -960 558634 480
rect 559626 -960 559738 480
rect 560730 -960 560842 480
rect 561834 -960 561946 480
<< via2 >>
rect 3422 694864 3478 694920
rect 3422 678136 3478 678192
rect 3422 661408 3478 661464
rect 3238 644680 3294 644736
rect 3422 627972 3478 628008
rect 3422 627952 3424 627972
rect 3424 627952 3476 627972
rect 3476 627952 3478 627972
rect 3422 611224 3478 611280
rect 3422 594496 3478 594552
rect 3054 577768 3110 577824
rect 3054 561040 3110 561096
rect 3330 510856 3386 510912
rect 3330 494128 3386 494184
rect 3146 477400 3202 477456
rect 3146 460672 3202 460728
rect 3330 443944 3386 444000
rect 3330 427216 3386 427272
rect 3330 410488 3386 410544
rect 3330 377032 3386 377088
rect 3330 360304 3386 360360
rect 3330 343576 3386 343632
rect 3330 326848 3386 326904
rect 3330 310120 3386 310176
rect 3330 293392 3386 293448
rect 3330 276664 3386 276720
rect 2962 259936 3018 259992
rect 3330 243208 3386 243264
rect 3330 226480 3386 226536
rect 3330 209788 3332 209808
rect 3332 209788 3384 209808
rect 3384 209788 3386 209808
rect 3330 209752 3386 209788
rect 3330 193024 3386 193080
rect 3054 176296 3110 176352
rect 3146 159568 3202 159624
rect 3514 544312 3570 544368
rect 3606 527584 3662 527640
rect 3606 393760 3662 393816
rect 3422 142840 3478 142896
rect 3330 126112 3386 126168
rect 2778 109384 2834 109440
rect 3882 92656 3938 92712
rect 3790 75928 3846 75984
rect 3698 59200 3754 59256
rect 3606 42472 3662 42528
rect 3514 25744 3570 25800
rect 3422 9016 3478 9072
rect 42982 7520 43038 7576
rect 46294 4800 46350 4856
rect 59358 87488 59414 87544
rect 59542 4936 59598 4992
rect 81530 104352 81586 104408
rect 81806 104352 81862 104408
rect 86866 152496 86922 152552
rect 85486 150456 85542 150512
rect 88062 152360 88118 152416
rect 97998 152088 98054 152144
rect 102690 152224 102746 152280
rect 105726 151816 105782 151872
rect 106830 151952 106886 152008
rect 110326 152632 110382 152688
rect 112626 151952 112682 152008
rect 119158 151816 119214 151872
rect 580170 695952 580226 696008
rect 580170 680348 580172 680368
rect 580172 680348 580224 680368
rect 580224 680348 580226 680368
rect 580170 680312 580226 680348
rect 580170 664672 580226 664728
rect 580170 649032 580226 649088
rect 580170 633428 580172 633448
rect 580172 633428 580224 633448
rect 580224 633428 580226 633448
rect 580170 633392 580226 633428
rect 580170 617752 580226 617808
rect 580170 602112 580226 602168
rect 580906 586508 580908 586528
rect 580908 586508 580960 586528
rect 580960 586508 580962 586528
rect 580906 586472 580962 586508
rect 580170 570832 580226 570888
rect 580170 555192 580226 555248
rect 580170 539588 580172 539608
rect 580172 539588 580224 539608
rect 580224 539588 580226 539608
rect 580170 539552 580226 539588
rect 580170 523912 580226 523968
rect 580170 508272 580226 508328
rect 580170 492668 580172 492688
rect 580172 492668 580224 492688
rect 580224 492668 580226 492688
rect 580170 492632 580226 492668
rect 580170 476992 580226 477048
rect 580170 461352 580226 461408
rect 580170 445748 580172 445768
rect 580172 445748 580224 445768
rect 580224 445748 580226 445768
rect 580170 445712 580226 445748
rect 580170 430072 580226 430128
rect 580170 414432 580226 414488
rect 580170 398828 580172 398848
rect 580172 398828 580224 398848
rect 580224 398828 580226 398848
rect 580170 398792 580226 398828
rect 580170 383152 580226 383208
rect 580170 367512 580226 367568
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 336232 580226 336288
rect 580170 320592 580226 320648
rect 580170 304988 580172 305008
rect 580172 304988 580224 305008
rect 580224 304988 580226 305008
rect 580170 304952 580226 304988
rect 580170 289312 580226 289368
rect 580170 273672 580226 273728
rect 580906 258068 580908 258088
rect 580908 258068 580960 258088
rect 580960 258068 580962 258088
rect 580906 258032 580962 258068
rect 580170 242392 580226 242448
rect 580170 226752 580226 226808
rect 580170 211148 580172 211168
rect 580172 211148 580224 211168
rect 580224 211148 580226 211168
rect 580170 211112 580226 211148
rect 580170 195472 580226 195528
rect 580170 179832 580226 179888
rect 580170 164228 580172 164248
rect 580172 164228 580224 164248
rect 580224 164228 580226 164248
rect 580170 164192 580226 164228
rect 124770 152088 124826 152144
rect 87510 149504 87566 149560
rect 94134 149504 94190 149560
rect 88062 149368 88118 149424
rect 83692 99864 83748 99920
rect 84428 99864 84484 99920
rect 83462 99332 83518 99388
rect 84290 99728 84346 99784
rect 84198 98232 84254 98288
rect 84888 99728 84944 99784
rect 85072 99864 85128 99920
rect 85532 99864 85588 99920
rect 85716 99864 85772 99920
rect 86360 99864 86416 99920
rect 86820 99864 86876 99920
rect 85210 99320 85266 99376
rect 85762 99728 85818 99784
rect 85670 98232 85726 98288
rect 85946 99592 86002 99648
rect 86314 99764 86316 99784
rect 86316 99764 86368 99784
rect 86368 99764 86370 99784
rect 86314 99728 86370 99764
rect 86498 98232 86554 98288
rect 86866 99592 86922 99648
rect 87464 99864 87520 99920
rect 87418 99592 87474 99648
rect 87326 99456 87382 99512
rect 88108 99864 88164 99920
rect 88062 99728 88118 99784
rect 88384 99762 88440 99818
rect 89120 99898 89176 99954
rect 87786 99456 87842 99512
rect 88062 99592 88118 99648
rect 88154 99456 88210 99512
rect 88522 99456 88578 99512
rect 89350 99592 89406 99648
rect 89856 99898 89912 99954
rect 90040 99864 90096 99920
rect 90684 99864 90740 99920
rect 89810 99592 89866 99648
rect 89626 97960 89682 98016
rect 89626 97824 89682 97880
rect 89902 98368 89958 98424
rect 90178 98232 90234 98288
rect 90362 99592 90418 99648
rect 90776 99728 90832 99784
rect 90730 99592 90786 99648
rect 90960 99898 91016 99954
rect 91190 99728 91246 99784
rect 91880 99898 91936 99954
rect 91834 99728 91890 99784
rect 91374 99592 91430 99648
rect 92248 99898 92304 99954
rect 92616 99898 92672 99954
rect 92800 99830 92856 99886
rect 92570 99592 92626 99648
rect 92202 98096 92258 98152
rect 92294 97960 92350 98016
rect 92754 99592 92810 99648
rect 93444 99728 93500 99784
rect 93628 99898 93684 99954
rect 93306 99592 93362 99648
rect 93122 97552 93178 97608
rect 93674 99592 93730 99648
rect 93398 98232 93454 98288
rect 94824 99864 94880 99920
rect 94042 99592 94098 99648
rect 94686 99764 94688 99784
rect 94688 99764 94740 99784
rect 94740 99764 94742 99784
rect 94686 99728 94742 99764
rect 95008 99728 95064 99784
rect 94502 88168 94558 88224
rect 95468 99864 95524 99920
rect 95652 99898 95708 99954
rect 95652 99728 95708 99784
rect 95146 97824 95202 97880
rect 95330 98232 95386 98288
rect 96204 99864 96260 99920
rect 96388 99728 96444 99784
rect 96756 99864 96812 99920
rect 97032 99898 97088 99954
rect 97216 99898 97272 99954
rect 97400 99898 97456 99954
rect 96618 99592 96674 99648
rect 96526 97552 96582 97608
rect 96986 99592 97042 99648
rect 97354 99728 97410 99784
rect 97538 99728 97594 99784
rect 98044 99898 98100 99954
rect 98320 99898 98376 99954
rect 98504 99898 98560 99954
rect 98780 99864 98836 99920
rect 97354 99592 97410 99648
rect 97538 97552 97594 97608
rect 97630 97416 97686 97472
rect 98274 99592 98330 99648
rect 97906 99492 97908 99512
rect 97908 99492 97960 99512
rect 97960 99492 97962 99512
rect 97906 99456 97962 99492
rect 97814 97144 97870 97200
rect 97538 96328 97594 96384
rect 98182 97552 98238 97608
rect 98090 97008 98146 97064
rect 98642 99592 98698 99648
rect 98642 97688 98698 97744
rect 98826 99456 98882 99512
rect 98918 97552 98974 97608
rect 99194 99728 99250 99784
rect 99700 99864 99756 99920
rect 99654 99764 99656 99784
rect 99656 99764 99708 99784
rect 99708 99764 99710 99784
rect 99102 97552 99158 97608
rect 99286 99592 99342 99648
rect 99010 97416 99066 97472
rect 98642 88984 98698 89040
rect 99654 99728 99710 99764
rect 99976 99864 100032 99920
rect 100344 99864 100400 99920
rect 100114 99592 100170 99648
rect 100206 98232 100262 98288
rect 100988 99898 101044 99954
rect 100666 98368 100722 98424
rect 100574 98096 100630 98152
rect 101632 99898 101688 99954
rect 101816 99898 101872 99954
rect 102000 99898 102056 99954
rect 102552 99898 102608 99954
rect 102736 99898 102792 99954
rect 103104 99898 103160 99954
rect 101402 99456 101458 99512
rect 101678 99592 101734 99648
rect 101954 99592 102010 99648
rect 101770 98232 101826 98288
rect 101770 95648 101826 95704
rect 102506 99728 102562 99784
rect 102874 99728 102930 99784
rect 102046 98232 102102 98288
rect 102046 95512 102102 95568
rect 102322 99456 102378 99512
rect 102782 99592 102838 99648
rect 103564 99864 103620 99920
rect 104208 99830 104264 99886
rect 103288 99764 103290 99784
rect 103290 99764 103342 99784
rect 103342 99764 103344 99784
rect 103288 99728 103344 99764
rect 104576 99864 104632 99920
rect 104944 99898 105000 99954
rect 103334 99628 103336 99648
rect 103336 99628 103388 99648
rect 103388 99628 103390 99648
rect 103334 99592 103390 99628
rect 103518 99592 103574 99648
rect 103058 98232 103114 98288
rect 103058 95512 103114 95568
rect 103150 91704 103206 91760
rect 103610 98232 103666 98288
rect 104162 99592 104218 99648
rect 104254 96464 104310 96520
rect 104530 99592 104586 99648
rect 104438 95648 104494 95704
rect 104070 95512 104126 95568
rect 104990 99728 105046 99784
rect 104622 95512 104678 95568
rect 104806 99628 104808 99648
rect 104808 99628 104860 99648
rect 104860 99628 104862 99648
rect 104806 99592 104862 99628
rect 104714 94424 104770 94480
rect 104438 87488 104494 87544
rect 105588 99864 105644 99920
rect 105266 98232 105322 98288
rect 106048 99898 106104 99954
rect 106094 96192 106150 96248
rect 106462 96600 106518 96656
rect 106738 96736 106794 96792
rect 107382 99864 107438 99920
rect 107520 99864 107576 99920
rect 107566 99728 107622 99784
rect 107888 99898 107944 99954
rect 107474 99592 107530 99648
rect 107290 96328 107346 96384
rect 107474 99456 107530 99512
rect 107658 99456 107714 99512
rect 107566 96192 107622 96248
rect 108256 99898 108312 99954
rect 108624 99898 108680 99954
rect 108394 99728 108450 99784
rect 107750 95376 107806 95432
rect 108808 99830 108864 99886
rect 109452 99864 109508 99920
rect 108302 99592 108358 99648
rect 108670 99592 108726 99648
rect 108762 99456 108818 99512
rect 108762 96600 108818 96656
rect 108670 96192 108726 96248
rect 110188 99864 110244 99920
rect 110648 99728 110704 99784
rect 110050 96192 110106 96248
rect 110326 98096 110382 98152
rect 110234 96736 110290 96792
rect 110602 99592 110658 99648
rect 110418 96464 110474 96520
rect 110142 93336 110198 93392
rect 111200 99864 111256 99920
rect 111384 99898 111440 99954
rect 111752 99864 111808 99920
rect 111706 99728 111762 99784
rect 111338 99456 111394 99512
rect 111614 99320 111670 99376
rect 111706 96328 111762 96384
rect 111430 95512 111486 95568
rect 105910 3440 105966 3496
rect 112074 99592 112130 99648
rect 112258 99320 112314 99376
rect 113316 99864 113372 99920
rect 112810 96872 112866 96928
rect 112718 96736 112774 96792
rect 112994 97008 113050 97064
rect 112902 96600 112958 96656
rect 113914 99456 113970 99512
rect 113914 97552 113970 97608
rect 114006 96600 114062 96656
rect 114328 99728 114384 99784
rect 114512 99864 114568 99920
rect 114190 96736 114246 96792
rect 114374 96872 114430 96928
rect 114374 96736 114430 96792
rect 114650 99592 114706 99648
rect 115018 99694 115074 99750
rect 115202 99332 115258 99388
rect 116168 99898 116224 99954
rect 116352 99898 116408 99954
rect 116536 99864 116592 99920
rect 116398 99728 116454 99784
rect 117088 99898 117144 99954
rect 115662 96736 115718 96792
rect 115570 96600 115626 96656
rect 116122 99456 116178 99512
rect 116766 97416 116822 97472
rect 118284 99864 118340 99920
rect 118468 99898 118524 99954
rect 118238 99748 118294 99784
rect 118238 99728 118240 99748
rect 118240 99728 118292 99748
rect 118292 99728 118294 99748
rect 117226 99592 117282 99648
rect 117226 99476 117282 99512
rect 117226 99456 117228 99476
rect 117228 99456 117280 99476
rect 117280 99456 117282 99476
rect 118928 99898 118984 99954
rect 118238 97008 118294 97064
rect 118698 99592 118754 99648
rect 118422 97144 118478 97200
rect 118330 96872 118386 96928
rect 119756 99864 119812 99920
rect 119618 99764 119620 99784
rect 119620 99764 119672 99784
rect 119672 99764 119674 99784
rect 119618 99728 119674 99764
rect 120078 99728 120134 99784
rect 120400 99898 120456 99954
rect 120768 99898 120824 99954
rect 121044 99898 121100 99954
rect 121504 99898 121560 99954
rect 121688 99830 121744 99886
rect 119802 97144 119858 97200
rect 119894 96056 119950 96112
rect 120446 99456 120502 99512
rect 122056 99864 122112 99920
rect 120998 97280 121054 97336
rect 121090 97144 121146 97200
rect 120630 96872 120686 96928
rect 121182 96872 121238 96928
rect 121642 99592 121698 99648
rect 121550 95920 121606 95976
rect 122516 99864 122572 99920
rect 122424 99728 122480 99784
rect 122194 99592 122250 99648
rect 122102 99456 122158 99512
rect 122562 98368 122618 98424
rect 122654 96736 122710 96792
rect 122470 4800 122526 4856
rect 123896 99864 123952 99920
rect 124264 99864 124320 99920
rect 124632 99864 124688 99920
rect 124034 98232 124090 98288
rect 123942 97552 123998 97608
rect 124402 99592 124458 99648
rect 125276 99864 125332 99920
rect 125230 96736 125286 96792
rect 125644 99898 125700 99954
rect 125920 99898 125976 99954
rect 126196 99898 126252 99954
rect 126472 99898 126528 99954
rect 125874 99592 125930 99648
rect 126656 99898 126712 99954
rect 125506 99456 125562 99512
rect 125782 99456 125838 99512
rect 125414 97008 125470 97064
rect 125046 92384 125102 92440
rect 125322 96600 125378 96656
rect 125598 99320 125654 99376
rect 126242 99592 126298 99648
rect 126150 99184 126206 99240
rect 126058 98232 126114 98288
rect 126886 98232 126942 98288
rect 126702 98096 126758 98152
rect 126610 97280 126666 97336
rect 124678 3304 124734 3360
rect 136086 152496 136142 152552
rect 129830 151816 129886 151872
rect 138662 152360 138718 152416
rect 580170 148552 580226 148608
rect 579986 132912 580042 132968
rect 580170 117272 580226 117328
rect 153198 94696 153254 94752
rect 140778 40840 140834 40896
rect 139398 18944 139454 19000
rect 157338 42064 157394 42120
rect 153290 28464 153346 28520
rect 156694 11736 156750 11792
rect 169850 40704 169906 40760
rect 173898 36352 173954 36408
rect 172518 20032 172574 20088
rect 190458 40568 190514 40624
rect 186318 37168 186374 37224
rect 189814 7520 189870 7576
rect 207018 38256 207074 38312
rect 202878 37032 202934 37088
rect 203062 9424 203118 9480
rect 206374 9288 206430 9344
rect 235998 94560 236054 94616
rect 223578 38120 223634 38176
rect 219438 24384 219494 24440
rect 219530 21392 219586 21448
rect 222934 6568 222990 6624
rect 240138 27104 240194 27160
rect 236182 9152 236238 9208
rect 239494 9016 239550 9072
rect 255318 25472 255374 25528
rect 256698 22888 256754 22944
rect 254950 8880 255006 8936
rect 270498 84904 270554 84960
rect 269118 26968 269174 27024
rect 273258 26832 273314 26888
rect 272614 10376 272670 10432
rect 289818 94424 289874 94480
rect 285770 28328 285826 28384
rect 285678 28192 285734 28248
rect 289174 10240 289230 10296
rect 335358 93472 335414 93528
rect 304998 84768 305054 84824
rect 306378 29552 306434 29608
rect 318798 31048 318854 31104
rect 322938 30912 322994 30968
rect 322294 13232 322350 13288
rect 321190 11600 321246 11656
rect 336738 39344 336794 39400
rect 339498 24248 339554 24304
rect 338854 13096 338910 13152
rect 356058 93336 356114 93392
rect 351918 24112 351974 24168
rect 368478 93200 368534 93256
rect 354310 12960 354366 13016
rect 372618 36896 372674 36952
rect 370870 14864 370926 14920
rect 371974 14728 372030 14784
rect 389178 93064 389234 93120
rect 385038 36760 385094 36816
rect 387430 14592 387486 14648
rect 388534 14456 388590 14512
rect 420918 90752 420974 90808
rect 405738 33768 405794 33824
rect 401690 32544 401746 32600
rect 403990 16088 404046 16144
rect 405094 15952 405150 16008
rect 436098 90616 436154 90672
rect 420550 15816 420606 15872
rect 434810 35672 434866 35728
rect 438858 37984 438914 38040
rect 437478 35536 437534 35592
rect 471978 96056 472034 96112
rect 451278 37848 451334 37904
rect 449898 17448 449954 17504
rect 451370 35400 451426 35456
rect 454038 35264 454094 35320
rect 452658 17312 452714 17368
rect 467930 32408 467986 32464
rect 470598 18808 470654 18864
rect 488538 95920 488594 95976
rect 485778 90480 485834 90536
rect 484398 35128 484454 35184
rect 484582 6432 484638 6488
rect 487894 6296 487950 6352
rect 502338 90344 502394 90400
rect 501050 17176 501106 17232
rect 505098 18672 505154 18728
rect 504454 6160 504510 6216
rect 521658 95784 521714 95840
rect 520278 21256 520334 21312
rect 519910 4800 519966 4856
rect 535458 79328 535514 79384
rect 534078 18536 534134 18592
rect 538218 36624 538274 36680
rect 536838 22752 536894 22808
rect 579618 70352 579674 70408
rect 552018 39208 552074 39264
rect 550730 19896 550786 19952
rect 554778 36488 554834 36544
rect 553398 22616 553454 22672
rect 580630 101632 580686 101688
rect 580538 85992 580594 86048
rect 580446 54712 580502 54768
rect 580354 23432 580410 23488
rect 580262 7792 580318 7848
<< metal3 >>
rect 580165 696010 580231 696013
rect 583520 696010 584960 696100
rect 580165 696008 584960 696010
rect 580165 695952 580170 696008
rect 580226 695952 584960 696008
rect 580165 695950 584960 695952
rect 580165 695947 580231 695950
rect 583520 695860 584960 695950
rect -960 694922 480 695012
rect 3417 694922 3483 694925
rect -960 694920 3483 694922
rect -960 694864 3422 694920
rect 3478 694864 3483 694920
rect -960 694862 3483 694864
rect -960 694772 480 694862
rect 3417 694859 3483 694862
rect 580165 680370 580231 680373
rect 583520 680370 584960 680460
rect 580165 680368 584960 680370
rect 580165 680312 580170 680368
rect 580226 680312 584960 680368
rect 580165 680310 584960 680312
rect 580165 680307 580231 680310
rect 583520 680220 584960 680310
rect -960 678194 480 678284
rect 3417 678194 3483 678197
rect -960 678192 3483 678194
rect -960 678136 3422 678192
rect 3478 678136 3483 678192
rect -960 678134 3483 678136
rect -960 678044 480 678134
rect 3417 678131 3483 678134
rect 580165 664730 580231 664733
rect 583520 664730 584960 664820
rect 580165 664728 584960 664730
rect 580165 664672 580170 664728
rect 580226 664672 584960 664728
rect 580165 664670 584960 664672
rect 580165 664667 580231 664670
rect 583520 664580 584960 664670
rect -960 661466 480 661556
rect 3417 661466 3483 661469
rect -960 661464 3483 661466
rect -960 661408 3422 661464
rect 3478 661408 3483 661464
rect -960 661406 3483 661408
rect -960 661316 480 661406
rect 3417 661403 3483 661406
rect 580165 649090 580231 649093
rect 583520 649090 584960 649180
rect 580165 649088 584960 649090
rect 580165 649032 580170 649088
rect 580226 649032 584960 649088
rect 580165 649030 584960 649032
rect 580165 649027 580231 649030
rect 583520 648940 584960 649030
rect -960 644738 480 644828
rect 3233 644738 3299 644741
rect -960 644736 3299 644738
rect -960 644680 3238 644736
rect 3294 644680 3299 644736
rect -960 644678 3299 644680
rect -960 644588 480 644678
rect 3233 644675 3299 644678
rect 580165 633450 580231 633453
rect 583520 633450 584960 633540
rect 580165 633448 584960 633450
rect 580165 633392 580170 633448
rect 580226 633392 584960 633448
rect 580165 633390 584960 633392
rect 580165 633387 580231 633390
rect 583520 633300 584960 633390
rect -960 628010 480 628100
rect 3417 628010 3483 628013
rect -960 628008 3483 628010
rect -960 627952 3422 628008
rect 3478 627952 3483 628008
rect -960 627950 3483 627952
rect -960 627860 480 627950
rect 3417 627947 3483 627950
rect 580165 617810 580231 617813
rect 583520 617810 584960 617900
rect 580165 617808 584960 617810
rect 580165 617752 580170 617808
rect 580226 617752 584960 617808
rect 580165 617750 584960 617752
rect 580165 617747 580231 617750
rect 583520 617660 584960 617750
rect -960 611282 480 611372
rect 3417 611282 3483 611285
rect -960 611280 3483 611282
rect -960 611224 3422 611280
rect 3478 611224 3483 611280
rect -960 611222 3483 611224
rect -960 611132 480 611222
rect 3417 611219 3483 611222
rect 580165 602170 580231 602173
rect 583520 602170 584960 602260
rect 580165 602168 584960 602170
rect 580165 602112 580170 602168
rect 580226 602112 584960 602168
rect 580165 602110 584960 602112
rect 580165 602107 580231 602110
rect 583520 602020 584960 602110
rect -960 594554 480 594644
rect 3417 594554 3483 594557
rect -960 594552 3483 594554
rect -960 594496 3422 594552
rect 3478 594496 3483 594552
rect -960 594494 3483 594496
rect -960 594404 480 594494
rect 3417 594491 3483 594494
rect 580901 586530 580967 586533
rect 583520 586530 584960 586620
rect 580901 586528 581010 586530
rect 580901 586472 580906 586528
rect 580962 586472 581010 586528
rect 580901 586467 581010 586472
rect 580950 586394 581010 586467
rect 582974 586470 584960 586530
rect 582974 586394 583034 586470
rect 580950 586334 583034 586394
rect 583520 586380 584960 586470
rect -960 577826 480 577916
rect 3049 577826 3115 577829
rect -960 577824 3115 577826
rect -960 577768 3054 577824
rect 3110 577768 3115 577824
rect -960 577766 3115 577768
rect -960 577676 480 577766
rect 3049 577763 3115 577766
rect 580165 570890 580231 570893
rect 583520 570890 584960 570980
rect 580165 570888 584960 570890
rect 580165 570832 580170 570888
rect 580226 570832 584960 570888
rect 580165 570830 584960 570832
rect 580165 570827 580231 570830
rect 583520 570740 584960 570830
rect -960 561098 480 561188
rect 3049 561098 3115 561101
rect -960 561096 3115 561098
rect -960 561040 3054 561096
rect 3110 561040 3115 561096
rect -960 561038 3115 561040
rect -960 560948 480 561038
rect 3049 561035 3115 561038
rect 580165 555250 580231 555253
rect 583520 555250 584960 555340
rect 580165 555248 584960 555250
rect 580165 555192 580170 555248
rect 580226 555192 584960 555248
rect 580165 555190 584960 555192
rect 580165 555187 580231 555190
rect 583520 555100 584960 555190
rect -960 544370 480 544460
rect 3509 544370 3575 544373
rect -960 544368 3575 544370
rect -960 544312 3514 544368
rect 3570 544312 3575 544368
rect -960 544310 3575 544312
rect -960 544220 480 544310
rect 3509 544307 3575 544310
rect 580165 539610 580231 539613
rect 583520 539610 584960 539700
rect 580165 539608 584960 539610
rect 580165 539552 580170 539608
rect 580226 539552 584960 539608
rect 580165 539550 584960 539552
rect 580165 539547 580231 539550
rect 583520 539460 584960 539550
rect -960 527642 480 527732
rect 3601 527642 3667 527645
rect -960 527640 3667 527642
rect -960 527584 3606 527640
rect 3662 527584 3667 527640
rect -960 527582 3667 527584
rect -960 527492 480 527582
rect 3601 527579 3667 527582
rect 580165 523970 580231 523973
rect 583520 523970 584960 524060
rect 580165 523968 584960 523970
rect 580165 523912 580170 523968
rect 580226 523912 584960 523968
rect 580165 523910 584960 523912
rect 580165 523907 580231 523910
rect 583520 523820 584960 523910
rect -960 510914 480 511004
rect 3325 510914 3391 510917
rect -960 510912 3391 510914
rect -960 510856 3330 510912
rect 3386 510856 3391 510912
rect -960 510854 3391 510856
rect -960 510764 480 510854
rect 3325 510851 3391 510854
rect 580165 508330 580231 508333
rect 583520 508330 584960 508420
rect 580165 508328 584960 508330
rect 580165 508272 580170 508328
rect 580226 508272 584960 508328
rect 580165 508270 584960 508272
rect 580165 508267 580231 508270
rect 583520 508180 584960 508270
rect -960 494186 480 494276
rect 3325 494186 3391 494189
rect -960 494184 3391 494186
rect -960 494128 3330 494184
rect 3386 494128 3391 494184
rect -960 494126 3391 494128
rect -960 494036 480 494126
rect 3325 494123 3391 494126
rect 580165 492690 580231 492693
rect 583520 492690 584960 492780
rect 580165 492688 584960 492690
rect 580165 492632 580170 492688
rect 580226 492632 584960 492688
rect 580165 492630 584960 492632
rect 580165 492627 580231 492630
rect 583520 492540 584960 492630
rect -960 477458 480 477548
rect 3141 477458 3207 477461
rect -960 477456 3207 477458
rect -960 477400 3146 477456
rect 3202 477400 3207 477456
rect -960 477398 3207 477400
rect -960 477308 480 477398
rect 3141 477395 3207 477398
rect 580165 477050 580231 477053
rect 583520 477050 584960 477140
rect 580165 477048 584960 477050
rect 580165 476992 580170 477048
rect 580226 476992 584960 477048
rect 580165 476990 584960 476992
rect 580165 476987 580231 476990
rect 583520 476900 584960 476990
rect 580165 461410 580231 461413
rect 583520 461410 584960 461500
rect 580165 461408 584960 461410
rect 580165 461352 580170 461408
rect 580226 461352 584960 461408
rect 580165 461350 584960 461352
rect 580165 461347 580231 461350
rect 583520 461260 584960 461350
rect -960 460730 480 460820
rect 3141 460730 3207 460733
rect -960 460728 3207 460730
rect -960 460672 3146 460728
rect 3202 460672 3207 460728
rect -960 460670 3207 460672
rect -960 460580 480 460670
rect 3141 460667 3207 460670
rect 580165 445770 580231 445773
rect 583520 445770 584960 445860
rect 580165 445768 584960 445770
rect 580165 445712 580170 445768
rect 580226 445712 584960 445768
rect 580165 445710 584960 445712
rect 580165 445707 580231 445710
rect 583520 445620 584960 445710
rect -960 444002 480 444092
rect 3325 444002 3391 444005
rect -960 444000 3391 444002
rect -960 443944 3330 444000
rect 3386 443944 3391 444000
rect -960 443942 3391 443944
rect -960 443852 480 443942
rect 3325 443939 3391 443942
rect 580165 430130 580231 430133
rect 583520 430130 584960 430220
rect 580165 430128 584960 430130
rect 580165 430072 580170 430128
rect 580226 430072 584960 430128
rect 580165 430070 584960 430072
rect 580165 430067 580231 430070
rect 583520 429980 584960 430070
rect -960 427274 480 427364
rect 3325 427274 3391 427277
rect -960 427272 3391 427274
rect -960 427216 3330 427272
rect 3386 427216 3391 427272
rect -960 427214 3391 427216
rect -960 427124 480 427214
rect 3325 427211 3391 427214
rect 580165 414490 580231 414493
rect 583520 414490 584960 414580
rect 580165 414488 584960 414490
rect 580165 414432 580170 414488
rect 580226 414432 584960 414488
rect 580165 414430 584960 414432
rect 580165 414427 580231 414430
rect 583520 414340 584960 414430
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 398850 580231 398853
rect 583520 398850 584960 398940
rect 580165 398848 584960 398850
rect 580165 398792 580170 398848
rect 580226 398792 584960 398848
rect 580165 398790 584960 398792
rect 580165 398787 580231 398790
rect 583520 398700 584960 398790
rect -960 393818 480 393908
rect 3601 393818 3667 393821
rect -960 393816 3667 393818
rect -960 393760 3606 393816
rect 3662 393760 3667 393816
rect -960 393758 3667 393760
rect -960 393668 480 393758
rect 3601 393755 3667 393758
rect 580165 383210 580231 383213
rect 583520 383210 584960 383300
rect 580165 383208 584960 383210
rect 580165 383152 580170 383208
rect 580226 383152 584960 383208
rect 580165 383150 584960 383152
rect 580165 383147 580231 383150
rect 583520 383060 584960 383150
rect -960 377090 480 377180
rect 3325 377090 3391 377093
rect -960 377088 3391 377090
rect -960 377032 3330 377088
rect 3386 377032 3391 377088
rect -960 377030 3391 377032
rect -960 376940 480 377030
rect 3325 377027 3391 377030
rect 580165 367570 580231 367573
rect 583520 367570 584960 367660
rect 580165 367568 584960 367570
rect 580165 367512 580170 367568
rect 580226 367512 584960 367568
rect 580165 367510 584960 367512
rect 580165 367507 580231 367510
rect 583520 367420 584960 367510
rect -960 360362 480 360452
rect 3325 360362 3391 360365
rect -960 360360 3391 360362
rect -960 360304 3330 360360
rect 3386 360304 3391 360360
rect -960 360302 3391 360304
rect -960 360212 480 360302
rect 3325 360299 3391 360302
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 343634 480 343724
rect 3325 343634 3391 343637
rect -960 343632 3391 343634
rect -960 343576 3330 343632
rect 3386 343576 3391 343632
rect -960 343574 3391 343576
rect -960 343484 480 343574
rect 3325 343571 3391 343574
rect 580165 336290 580231 336293
rect 583520 336290 584960 336380
rect 580165 336288 584960 336290
rect 580165 336232 580170 336288
rect 580226 336232 584960 336288
rect 580165 336230 584960 336232
rect 580165 336227 580231 336230
rect 583520 336140 584960 336230
rect -960 326906 480 326996
rect 3325 326906 3391 326909
rect -960 326904 3391 326906
rect -960 326848 3330 326904
rect 3386 326848 3391 326904
rect -960 326846 3391 326848
rect -960 326756 480 326846
rect 3325 326843 3391 326846
rect 580165 320650 580231 320653
rect 583520 320650 584960 320740
rect 580165 320648 584960 320650
rect 580165 320592 580170 320648
rect 580226 320592 584960 320648
rect 580165 320590 584960 320592
rect 580165 320587 580231 320590
rect 583520 320500 584960 320590
rect -960 310178 480 310268
rect 3325 310178 3391 310181
rect -960 310176 3391 310178
rect -960 310120 3330 310176
rect 3386 310120 3391 310176
rect -960 310118 3391 310120
rect -960 310028 480 310118
rect 3325 310115 3391 310118
rect 580165 305010 580231 305013
rect 583520 305010 584960 305100
rect 580165 305008 584960 305010
rect 580165 304952 580170 305008
rect 580226 304952 584960 305008
rect 580165 304950 584960 304952
rect 580165 304947 580231 304950
rect 583520 304860 584960 304950
rect -960 293450 480 293540
rect 3325 293450 3391 293453
rect -960 293448 3391 293450
rect -960 293392 3330 293448
rect 3386 293392 3391 293448
rect -960 293390 3391 293392
rect -960 293300 480 293390
rect 3325 293387 3391 293390
rect 580165 289370 580231 289373
rect 583520 289370 584960 289460
rect 580165 289368 584960 289370
rect 580165 289312 580170 289368
rect 580226 289312 584960 289368
rect 580165 289310 584960 289312
rect 580165 289307 580231 289310
rect 583520 289220 584960 289310
rect -960 276722 480 276812
rect 3325 276722 3391 276725
rect -960 276720 3391 276722
rect -960 276664 3330 276720
rect 3386 276664 3391 276720
rect -960 276662 3391 276664
rect -960 276572 480 276662
rect 3325 276659 3391 276662
rect 580165 273730 580231 273733
rect 583520 273730 584960 273820
rect 580165 273728 584960 273730
rect 580165 273672 580170 273728
rect 580226 273672 584960 273728
rect 580165 273670 584960 273672
rect 580165 273667 580231 273670
rect 583520 273580 584960 273670
rect -960 259994 480 260084
rect 2957 259994 3023 259997
rect -960 259992 3023 259994
rect -960 259936 2962 259992
rect 3018 259936 3023 259992
rect -960 259934 3023 259936
rect -960 259844 480 259934
rect 2957 259931 3023 259934
rect 580901 258090 580967 258093
rect 583520 258090 584960 258180
rect 580901 258088 581010 258090
rect 580901 258032 580906 258088
rect 580962 258032 581010 258088
rect 580901 258027 581010 258032
rect 580950 257954 581010 258027
rect 582974 258030 584960 258090
rect 582974 257954 583034 258030
rect 580950 257894 583034 257954
rect 583520 257940 584960 258030
rect -960 243266 480 243356
rect 3325 243266 3391 243269
rect -960 243264 3391 243266
rect -960 243208 3330 243264
rect 3386 243208 3391 243264
rect -960 243206 3391 243208
rect -960 243116 480 243206
rect 3325 243203 3391 243206
rect 580165 242450 580231 242453
rect 583520 242450 584960 242540
rect 580165 242448 584960 242450
rect 580165 242392 580170 242448
rect 580226 242392 584960 242448
rect 580165 242390 584960 242392
rect 580165 242387 580231 242390
rect 583520 242300 584960 242390
rect 580165 226810 580231 226813
rect 583520 226810 584960 226900
rect 580165 226808 584960 226810
rect 580165 226752 580170 226808
rect 580226 226752 584960 226808
rect 580165 226750 584960 226752
rect 580165 226747 580231 226750
rect 583520 226660 584960 226750
rect -960 226538 480 226628
rect 3325 226538 3391 226541
rect -960 226536 3391 226538
rect -960 226480 3330 226536
rect 3386 226480 3391 226536
rect -960 226478 3391 226480
rect -960 226388 480 226478
rect 3325 226475 3391 226478
rect 580165 211170 580231 211173
rect 583520 211170 584960 211260
rect 580165 211168 584960 211170
rect 580165 211112 580170 211168
rect 580226 211112 584960 211168
rect 580165 211110 584960 211112
rect 580165 211107 580231 211110
rect 583520 211020 584960 211110
rect -960 209810 480 209900
rect 3325 209810 3391 209813
rect -960 209808 3391 209810
rect -960 209752 3330 209808
rect 3386 209752 3391 209808
rect -960 209750 3391 209752
rect -960 209660 480 209750
rect 3325 209747 3391 209750
rect 580165 195530 580231 195533
rect 583520 195530 584960 195620
rect 580165 195528 584960 195530
rect 580165 195472 580170 195528
rect 580226 195472 584960 195528
rect 580165 195470 584960 195472
rect 580165 195467 580231 195470
rect 583520 195380 584960 195470
rect -960 193082 480 193172
rect 3325 193082 3391 193085
rect -960 193080 3391 193082
rect -960 193024 3330 193080
rect 3386 193024 3391 193080
rect -960 193022 3391 193024
rect -960 192932 480 193022
rect 3325 193019 3391 193022
rect 580165 179890 580231 179893
rect 583520 179890 584960 179980
rect 580165 179888 584960 179890
rect 580165 179832 580170 179888
rect 580226 179832 584960 179888
rect 580165 179830 584960 179832
rect 580165 179827 580231 179830
rect 583520 179740 584960 179830
rect -960 176354 480 176444
rect 3049 176354 3115 176357
rect -960 176352 3115 176354
rect -960 176296 3054 176352
rect 3110 176296 3115 176352
rect -960 176294 3115 176296
rect -960 176204 480 176294
rect 3049 176291 3115 176294
rect 580165 164250 580231 164253
rect 583520 164250 584960 164340
rect 580165 164248 584960 164250
rect 580165 164192 580170 164248
rect 580226 164192 584960 164248
rect 580165 164190 584960 164192
rect 580165 164187 580231 164190
rect 583520 164100 584960 164190
rect -960 159626 480 159716
rect 3141 159626 3207 159629
rect -960 159624 3207 159626
rect -960 159568 3146 159624
rect 3202 159568 3207 159624
rect -960 159566 3207 159568
rect -960 159476 480 159566
rect 3141 159563 3207 159566
rect 110321 152690 110387 152693
rect 122598 152690 122604 152692
rect 110321 152688 122604 152690
rect 110321 152632 110326 152688
rect 110382 152632 122604 152688
rect 110321 152630 122604 152632
rect 110321 152627 110387 152630
rect 122598 152628 122604 152630
rect 122668 152628 122674 152692
rect 86861 152554 86927 152557
rect 136081 152554 136147 152557
rect 86861 152552 136147 152554
rect 86861 152496 86866 152552
rect 86922 152496 136086 152552
rect 136142 152496 136147 152552
rect 86861 152494 136147 152496
rect 86861 152491 86927 152494
rect 136081 152491 136147 152494
rect 88057 152418 88123 152421
rect 138657 152418 138723 152421
rect 88057 152416 138723 152418
rect 88057 152360 88062 152416
rect 88118 152360 138662 152416
rect 138718 152360 138723 152416
rect 88057 152358 138723 152360
rect 88057 152355 88123 152358
rect 138657 152355 138723 152358
rect 102685 152282 102751 152285
rect 124254 152282 124260 152284
rect 102685 152280 124260 152282
rect 102685 152224 102690 152280
rect 102746 152224 124260 152280
rect 102685 152222 124260 152224
rect 102685 152219 102751 152222
rect 124254 152220 124260 152222
rect 124324 152220 124330 152284
rect 97993 152146 98059 152149
rect 124765 152146 124831 152149
rect 97993 152144 124831 152146
rect 97993 152088 97998 152144
rect 98054 152088 124770 152144
rect 124826 152088 124831 152144
rect 97993 152086 124831 152088
rect 97993 152083 98059 152086
rect 124765 152083 124831 152086
rect 83774 151948 83780 152012
rect 83844 152010 83850 152012
rect 106825 152010 106891 152013
rect 83844 152008 106891 152010
rect 83844 151952 106830 152008
rect 106886 151952 106891 152008
rect 83844 151950 106891 151952
rect 83844 151948 83850 151950
rect 106825 151947 106891 151950
rect 112621 152010 112687 152013
rect 124438 152010 124444 152012
rect 112621 152008 124444 152010
rect 112621 151952 112626 152008
rect 112682 151952 124444 152008
rect 112621 151950 124444 151952
rect 112621 151947 112687 151950
rect 124438 151948 124444 151950
rect 124508 151948 124514 152012
rect 82486 151812 82492 151876
rect 82556 151874 82562 151876
rect 105721 151874 105787 151877
rect 82556 151872 105787 151874
rect 82556 151816 105726 151872
rect 105782 151816 105787 151872
rect 82556 151814 105787 151816
rect 82556 151812 82562 151814
rect 105721 151811 105787 151814
rect 119153 151874 119219 151877
rect 129825 151874 129891 151877
rect 119153 151872 129891 151874
rect 119153 151816 119158 151872
rect 119214 151816 129830 151872
rect 129886 151816 129891 151872
rect 119153 151814 129891 151816
rect 119153 151811 119219 151814
rect 129825 151811 129891 151814
rect 85481 150514 85547 150517
rect 128854 150514 128860 150516
rect 85481 150512 128860 150514
rect 85481 150456 85486 150512
rect 85542 150456 128860 150512
rect 85481 150454 128860 150456
rect 85481 150451 85547 150454
rect 128854 150452 128860 150454
rect 128924 150452 128930 150516
rect 87505 149562 87571 149565
rect 94129 149562 94195 149565
rect 87505 149560 94195 149562
rect 87505 149504 87510 149560
rect 87566 149504 94134 149560
rect 94190 149504 94195 149560
rect 87505 149502 94195 149504
rect 87505 149499 87571 149502
rect 94129 149499 94195 149502
rect 83958 149364 83964 149428
rect 84028 149426 84034 149428
rect 88057 149426 88123 149429
rect 84028 149424 88123 149426
rect 84028 149368 88062 149424
rect 88118 149368 88123 149424
rect 84028 149366 88123 149368
rect 84028 149364 84034 149366
rect 88057 149363 88123 149366
rect 580165 148610 580231 148613
rect 583520 148610 584960 148700
rect 580165 148608 584960 148610
rect 580165 148552 580170 148608
rect 580226 148552 584960 148608
rect 580165 148550 584960 148552
rect 580165 148547 580231 148550
rect 583520 148460 584960 148550
rect -960 142898 480 142988
rect 3417 142898 3483 142901
rect -960 142896 3483 142898
rect -960 142840 3422 142896
rect 3478 142840 3483 142896
rect -960 142838 3483 142840
rect -960 142748 480 142838
rect 3417 142835 3483 142838
rect 579981 132970 580047 132973
rect 583520 132970 584960 133060
rect 579981 132968 584960 132970
rect 579981 132912 579986 132968
rect 580042 132912 584960 132968
rect 579981 132910 584960 132912
rect 579981 132907 580047 132910
rect 583520 132820 584960 132910
rect -960 126170 480 126260
rect 3325 126170 3391 126173
rect -960 126168 3391 126170
rect -960 126112 3330 126168
rect 3386 126112 3391 126168
rect -960 126110 3391 126112
rect -960 126020 480 126110
rect 3325 126107 3391 126110
rect 580165 117330 580231 117333
rect 583520 117330 584960 117420
rect 580165 117328 584960 117330
rect 580165 117272 580170 117328
rect 580226 117272 584960 117328
rect 580165 117270 584960 117272
rect 580165 117267 580231 117270
rect 583520 117180 584960 117270
rect -960 109442 480 109532
rect 2773 109442 2839 109445
rect -960 109440 2839 109442
rect -960 109384 2778 109440
rect 2834 109384 2839 109440
rect -960 109382 2839 109384
rect -960 109292 480 109382
rect 2773 109379 2839 109382
rect 81525 104410 81591 104413
rect 81801 104410 81867 104413
rect 81525 104408 81867 104410
rect 81525 104352 81530 104408
rect 81586 104352 81806 104408
rect 81862 104352 81867 104408
rect 81525 104350 81867 104352
rect 81525 104347 81591 104350
rect 81801 104347 81867 104350
rect 580625 101690 580691 101693
rect 583520 101690 584960 101780
rect 580625 101688 584960 101690
rect 580625 101632 580630 101688
rect 580686 101632 584960 101688
rect 580625 101630 584960 101632
rect 580625 101627 580691 101630
rect 583520 101540 584960 101630
rect 99782 100132 99788 100196
rect 99852 100194 99858 100196
rect 124438 100194 124444 100196
rect 99852 100134 111810 100194
rect 99852 100132 99858 100134
rect 83774 99996 83780 100060
rect 83844 100058 83850 100060
rect 110638 100058 110644 100060
rect 83844 99998 88810 100058
rect 83844 99996 83850 99998
rect 83687 99922 83753 99925
rect 83414 99920 83753 99922
rect 83414 99864 83692 99920
rect 83748 99864 83753 99920
rect 83414 99862 83753 99864
rect 83414 99393 83474 99862
rect 83687 99859 83753 99862
rect 84142 99860 84148 99924
rect 84212 99922 84218 99924
rect 84423 99922 84489 99925
rect 85067 99924 85133 99925
rect 85062 99922 85068 99924
rect 84212 99920 84489 99922
rect 84212 99864 84428 99920
rect 84484 99864 84489 99920
rect 84212 99862 84489 99864
rect 84976 99862 85068 99922
rect 84212 99860 84218 99862
rect 84423 99859 84489 99862
rect 85062 99860 85068 99862
rect 85132 99860 85138 99924
rect 85527 99922 85593 99925
rect 85711 99922 85777 99925
rect 86355 99924 86421 99925
rect 86350 99922 86356 99924
rect 85527 99920 85636 99922
rect 85527 99864 85532 99920
rect 85588 99864 85636 99920
rect 85067 99859 85133 99860
rect 85527 99859 85636 99864
rect 85711 99920 86004 99922
rect 85711 99864 85716 99920
rect 85772 99864 86004 99920
rect 85711 99862 86004 99864
rect 86264 99862 86356 99922
rect 85711 99859 85777 99862
rect 84285 99786 84351 99789
rect 84883 99786 84949 99789
rect 84285 99784 84949 99786
rect 84285 99728 84290 99784
rect 84346 99728 84888 99784
rect 84944 99728 84949 99784
rect 84285 99726 84949 99728
rect 85576 99788 85636 99859
rect 85576 99726 85620 99788
rect 84285 99723 84351 99726
rect 84883 99723 84949 99726
rect 85614 99724 85620 99726
rect 85684 99724 85690 99788
rect 85757 99786 85823 99789
rect 85944 99786 86004 99862
rect 86350 99860 86356 99862
rect 86420 99860 86426 99924
rect 86815 99922 86881 99925
rect 87459 99922 87525 99925
rect 88103 99922 88169 99925
rect 86542 99920 86881 99922
rect 86542 99864 86820 99920
rect 86876 99864 86881 99920
rect 86542 99862 86881 99864
rect 86355 99859 86421 99860
rect 86309 99786 86375 99789
rect 85757 99784 86004 99786
rect 85757 99728 85762 99784
rect 85818 99728 86004 99784
rect 85757 99726 86004 99728
rect 86174 99784 86375 99786
rect 86174 99728 86314 99784
rect 86370 99728 86375 99784
rect 86174 99726 86375 99728
rect 85757 99723 85823 99726
rect 85941 99650 86007 99653
rect 86174 99650 86234 99726
rect 86309 99723 86375 99726
rect 85941 99648 86234 99650
rect 85941 99592 85946 99648
rect 86002 99592 86234 99648
rect 85941 99590 86234 99592
rect 86542 99650 86602 99862
rect 86815 99859 86881 99862
rect 87278 99920 87525 99922
rect 87278 99864 87464 99920
rect 87520 99864 87525 99920
rect 87278 99862 87525 99864
rect 86861 99650 86927 99653
rect 86542 99648 86927 99650
rect 86542 99592 86866 99648
rect 86922 99592 86927 99648
rect 86542 99590 86927 99592
rect 85941 99587 86007 99590
rect 86861 99587 86927 99590
rect 87278 99517 87338 99862
rect 87459 99859 87525 99862
rect 87922 99920 88169 99922
rect 87922 99864 88108 99920
rect 88164 99864 88169 99920
rect 87922 99862 88169 99864
rect 87413 99650 87479 99653
rect 87922 99650 87982 99862
rect 88103 99859 88169 99862
rect 88379 99818 88445 99823
rect 88057 99786 88123 99789
rect 88057 99784 88258 99786
rect 88057 99728 88062 99784
rect 88118 99728 88258 99784
rect 88379 99762 88384 99818
rect 88440 99762 88445 99818
rect 88379 99757 88445 99762
rect 88057 99726 88258 99728
rect 88057 99723 88123 99726
rect 88057 99650 88123 99653
rect 87413 99648 87844 99650
rect 87413 99592 87418 99648
rect 87474 99592 87844 99648
rect 87413 99590 87844 99592
rect 87922 99648 88123 99650
rect 87922 99592 88062 99648
rect 88118 99592 88123 99648
rect 87922 99590 88123 99592
rect 87413 99587 87479 99590
rect 87784 99517 87844 99590
rect 88057 99587 88123 99590
rect 88198 99517 88258 99726
rect 87278 99512 87387 99517
rect 87278 99456 87326 99512
rect 87382 99456 87387 99512
rect 87278 99454 87387 99456
rect 87321 99451 87387 99454
rect 87781 99512 87847 99517
rect 87781 99456 87786 99512
rect 87842 99456 87847 99512
rect 87781 99451 87847 99456
rect 88149 99512 88258 99517
rect 88149 99456 88154 99512
rect 88210 99456 88258 99512
rect 88149 99454 88258 99456
rect 88382 99514 88442 99757
rect 88517 99514 88583 99517
rect 88382 99512 88583 99514
rect 88382 99456 88522 99512
rect 88578 99456 88583 99512
rect 88382 99454 88583 99456
rect 88750 99514 88810 99998
rect 108668 99998 109050 100058
rect 108668 99959 108728 99998
rect 89115 99954 89181 99959
rect 89115 99924 89120 99954
rect 89176 99924 89181 99954
rect 89851 99954 89917 99959
rect 89110 99860 89116 99924
rect 89180 99922 89186 99924
rect 89180 99862 89238 99922
rect 89851 99898 89856 99954
rect 89912 99898 89917 99954
rect 90955 99954 91021 99959
rect 90035 99924 90101 99925
rect 89851 99893 89917 99898
rect 89180 99860 89186 99862
rect 89854 99653 89914 99893
rect 90030 99860 90036 99924
rect 90100 99922 90106 99924
rect 90679 99922 90745 99925
rect 90955 99924 90960 99954
rect 91016 99924 91021 99954
rect 91875 99954 91941 99959
rect 90100 99862 90192 99922
rect 90406 99920 90745 99922
rect 90406 99864 90684 99920
rect 90740 99864 90745 99920
rect 90406 99862 90745 99864
rect 90100 99860 90106 99862
rect 90035 99859 90101 99860
rect 90406 99653 90466 99862
rect 90679 99859 90745 99862
rect 90950 99860 90956 99924
rect 91020 99922 91026 99924
rect 91020 99862 91078 99922
rect 91875 99898 91880 99954
rect 91936 99898 91941 99954
rect 91875 99893 91941 99898
rect 92243 99954 92309 99959
rect 92243 99898 92248 99954
rect 92304 99898 92309 99954
rect 92243 99893 92309 99898
rect 92611 99954 92677 99959
rect 92611 99898 92616 99954
rect 92672 99898 92677 99954
rect 93623 99954 93689 99959
rect 95647 99956 95713 99959
rect 92611 99893 92677 99898
rect 91020 99860 91026 99862
rect 91878 99789 91938 99893
rect 90771 99788 90837 99789
rect 90766 99786 90772 99788
rect 90680 99726 90772 99786
rect 90766 99724 90772 99726
rect 90836 99724 90842 99788
rect 91185 99786 91251 99789
rect 91142 99784 91251 99786
rect 91142 99728 91190 99784
rect 91246 99728 91251 99784
rect 90771 99723 90837 99724
rect 91142 99723 91251 99728
rect 91829 99784 91938 99789
rect 91829 99728 91834 99784
rect 91890 99728 91938 99784
rect 91829 99726 91938 99728
rect 91829 99723 91895 99726
rect 89345 99650 89411 99653
rect 89478 99650 89484 99652
rect 89345 99648 89484 99650
rect 89345 99592 89350 99648
rect 89406 99592 89484 99648
rect 89345 99590 89484 99592
rect 89345 99587 89411 99590
rect 89478 99588 89484 99590
rect 89548 99588 89554 99652
rect 89805 99648 89914 99653
rect 89805 99592 89810 99648
rect 89866 99592 89914 99648
rect 89805 99590 89914 99592
rect 90357 99648 90466 99653
rect 90357 99592 90362 99648
rect 90418 99592 90466 99648
rect 90357 99590 90466 99592
rect 89805 99587 89871 99590
rect 90357 99587 90423 99590
rect 90582 99588 90588 99652
rect 90652 99650 90658 99652
rect 90725 99650 90791 99653
rect 90652 99648 90791 99650
rect 90652 99592 90730 99648
rect 90786 99592 90791 99648
rect 90652 99590 90791 99592
rect 91142 99650 91202 99723
rect 91369 99650 91435 99653
rect 91142 99648 91435 99650
rect 91142 99592 91374 99648
rect 91430 99592 91435 99648
rect 91142 99590 91435 99592
rect 90652 99588 90658 99590
rect 90725 99587 90791 99590
rect 91369 99587 91435 99590
rect 91502 99588 91508 99652
rect 91572 99650 91578 99652
rect 92246 99650 92306 99893
rect 92614 99653 92674 99893
rect 92795 99886 92861 99891
rect 92795 99830 92800 99886
rect 92856 99830 92861 99886
rect 93342 99860 93348 99924
rect 93412 99922 93418 99924
rect 93623 99922 93628 99954
rect 93412 99898 93628 99922
rect 93684 99898 93689 99954
rect 95604 99954 95713 99956
rect 93412 99893 93689 99898
rect 93412 99862 93686 99893
rect 93412 99860 93418 99862
rect 94446 99860 94452 99924
rect 94516 99922 94522 99924
rect 94819 99922 94885 99925
rect 94516 99920 94885 99922
rect 94516 99864 94824 99920
rect 94880 99864 94885 99920
rect 94516 99862 94885 99864
rect 94516 99860 94522 99862
rect 94819 99859 94885 99862
rect 95182 99860 95188 99924
rect 95252 99922 95258 99924
rect 95463 99922 95529 99925
rect 95252 99920 95529 99922
rect 95252 99864 95468 99920
rect 95524 99864 95529 99920
rect 95252 99862 95529 99864
rect 95252 99860 95258 99862
rect 95463 99859 95529 99862
rect 95604 99898 95652 99954
rect 95708 99898 95713 99954
rect 97027 99954 97093 99959
rect 95604 99893 95713 99898
rect 92795 99825 92861 99830
rect 92798 99653 92858 99825
rect 95604 99789 95664 99893
rect 95918 99860 95924 99924
rect 95988 99922 95994 99924
rect 96199 99922 96265 99925
rect 96751 99922 96817 99925
rect 95988 99920 96265 99922
rect 95988 99864 96204 99920
rect 96260 99864 96265 99920
rect 95988 99862 96265 99864
rect 95988 99860 95994 99862
rect 96199 99859 96265 99862
rect 96570 99920 96817 99922
rect 96570 99864 96756 99920
rect 96812 99864 96817 99920
rect 97027 99898 97032 99954
rect 97088 99898 97093 99954
rect 97027 99893 97093 99898
rect 97211 99954 97277 99959
rect 97211 99898 97216 99954
rect 97272 99898 97277 99954
rect 97211 99893 97277 99898
rect 97395 99954 97461 99959
rect 97395 99898 97400 99954
rect 97456 99898 97461 99954
rect 97395 99893 97461 99898
rect 98039 99956 98105 99959
rect 98039 99954 98148 99956
rect 98039 99898 98044 99954
rect 98100 99924 98148 99954
rect 98315 99954 98381 99959
rect 98100 99898 98132 99924
rect 98039 99893 98132 99898
rect 96570 99862 96817 99864
rect 93439 99786 93505 99789
rect 94681 99788 94747 99789
rect 95003 99788 95069 99789
rect 93710 99786 93716 99788
rect 93439 99784 93716 99786
rect 93439 99728 93444 99784
rect 93500 99728 93716 99784
rect 93439 99726 93716 99728
rect 93439 99723 93505 99726
rect 93710 99724 93716 99726
rect 93780 99724 93786 99788
rect 94630 99786 94636 99788
rect 94590 99726 94636 99786
rect 94700 99784 94747 99788
rect 94998 99786 95004 99788
rect 94742 99728 94747 99784
rect 94630 99724 94636 99726
rect 94700 99724 94747 99728
rect 94912 99726 95004 99786
rect 94998 99724 95004 99726
rect 95068 99724 95074 99788
rect 95604 99784 95713 99789
rect 95604 99728 95652 99784
rect 95708 99728 95713 99784
rect 95604 99726 95713 99728
rect 94681 99723 94747 99724
rect 95003 99723 95069 99724
rect 95647 99723 95713 99726
rect 96102 99724 96108 99788
rect 96172 99786 96178 99788
rect 96383 99786 96449 99789
rect 96172 99784 96449 99786
rect 96172 99728 96388 99784
rect 96444 99728 96449 99784
rect 96172 99726 96449 99728
rect 96172 99724 96178 99726
rect 96383 99723 96449 99726
rect 96570 99653 96630 99862
rect 96751 99859 96817 99862
rect 97030 99653 97090 99893
rect 91572 99590 92306 99650
rect 92565 99648 92674 99653
rect 92565 99592 92570 99648
rect 92626 99592 92674 99648
rect 92565 99590 92674 99592
rect 92749 99648 92858 99653
rect 92749 99592 92754 99648
rect 92810 99592 92858 99648
rect 92749 99590 92858 99592
rect 93301 99650 93367 99653
rect 93526 99650 93532 99652
rect 93301 99648 93532 99650
rect 93301 99592 93306 99648
rect 93362 99592 93532 99648
rect 93301 99590 93532 99592
rect 91572 99588 91578 99590
rect 92565 99587 92631 99590
rect 92749 99587 92815 99590
rect 93301 99587 93367 99590
rect 93526 99588 93532 99590
rect 93596 99588 93602 99652
rect 93669 99650 93735 99653
rect 94037 99650 94103 99653
rect 93669 99648 94103 99650
rect 93669 99592 93674 99648
rect 93730 99592 94042 99648
rect 94098 99592 94103 99648
rect 93669 99590 94103 99592
rect 96570 99648 96679 99653
rect 96570 99592 96618 99648
rect 96674 99592 96679 99648
rect 96570 99590 96679 99592
rect 93669 99587 93735 99590
rect 94037 99587 94103 99590
rect 96613 99587 96679 99590
rect 96981 99648 97090 99653
rect 96981 99592 96986 99648
rect 97042 99592 97090 99648
rect 96981 99590 97090 99592
rect 97214 99650 97274 99893
rect 97398 99789 97458 99893
rect 98088 99862 98132 99893
rect 98126 99860 98132 99862
rect 98196 99860 98202 99924
rect 98315 99898 98320 99954
rect 98376 99898 98381 99954
rect 98315 99893 98381 99898
rect 98499 99954 98565 99959
rect 98499 99898 98504 99954
rect 98560 99898 98565 99954
rect 100983 99956 101049 99959
rect 100983 99954 101092 99956
rect 98499 99893 98565 99898
rect 98775 99922 98841 99925
rect 99695 99922 99761 99925
rect 98775 99920 99252 99922
rect 97349 99784 97458 99789
rect 97349 99728 97354 99784
rect 97410 99728 97458 99784
rect 97349 99726 97458 99728
rect 97533 99786 97599 99789
rect 97758 99786 97764 99788
rect 97533 99784 97764 99786
rect 97533 99728 97538 99784
rect 97594 99728 97764 99784
rect 97533 99726 97764 99728
rect 97349 99723 97415 99726
rect 97533 99723 97599 99726
rect 97758 99724 97764 99726
rect 97828 99724 97834 99788
rect 98318 99653 98378 99893
rect 97349 99650 97415 99653
rect 97214 99648 97415 99650
rect 97214 99592 97354 99648
rect 97410 99592 97415 99648
rect 97214 99590 97415 99592
rect 96981 99587 97047 99590
rect 97349 99587 97415 99590
rect 98269 99648 98378 99653
rect 98269 99592 98274 99648
rect 98330 99592 98378 99648
rect 98269 99590 98378 99592
rect 98502 99650 98562 99893
rect 98775 99864 98780 99920
rect 98836 99864 99252 99920
rect 98775 99862 99252 99864
rect 98775 99859 98841 99862
rect 99192 99789 99252 99862
rect 99422 99920 99761 99922
rect 99422 99864 99700 99920
rect 99756 99864 99761 99920
rect 99422 99862 99761 99864
rect 99189 99784 99255 99789
rect 99189 99728 99194 99784
rect 99250 99728 99255 99784
rect 99189 99723 99255 99728
rect 98637 99650 98703 99653
rect 98502 99648 98703 99650
rect 98502 99592 98642 99648
rect 98698 99592 98703 99648
rect 98502 99590 98703 99592
rect 98269 99587 98335 99590
rect 98637 99587 98703 99590
rect 99281 99650 99347 99653
rect 99422 99650 99482 99862
rect 99695 99859 99761 99862
rect 99971 99920 100037 99925
rect 99971 99864 99976 99920
rect 100032 99864 100037 99920
rect 99971 99859 100037 99864
rect 100339 99922 100405 99925
rect 100518 99922 100524 99924
rect 100339 99920 100524 99922
rect 100339 99864 100344 99920
rect 100400 99864 100524 99920
rect 100339 99862 100524 99864
rect 100339 99859 100405 99862
rect 100518 99860 100524 99862
rect 100588 99860 100594 99924
rect 100983 99898 100988 99954
rect 101044 99898 101092 99954
rect 101627 99954 101693 99959
rect 101627 99922 101632 99954
rect 100983 99893 101092 99898
rect 99649 99786 99715 99789
rect 99782 99786 99788 99788
rect 99649 99784 99788 99786
rect 99649 99728 99654 99784
rect 99710 99728 99788 99784
rect 99649 99726 99788 99728
rect 99649 99723 99715 99726
rect 99782 99724 99788 99726
rect 99852 99724 99858 99788
rect 99281 99648 99482 99650
rect 99281 99592 99286 99648
rect 99342 99592 99482 99648
rect 99281 99590 99482 99592
rect 99974 99650 100034 99859
rect 100109 99650 100175 99653
rect 99974 99648 100175 99650
rect 99974 99592 100114 99648
rect 100170 99592 100175 99648
rect 99974 99590 100175 99592
rect 99281 99587 99347 99590
rect 100109 99587 100175 99590
rect 97901 99514 97967 99517
rect 88750 99512 97967 99514
rect 88750 99456 97906 99512
rect 97962 99456 97967 99512
rect 88750 99454 97967 99456
rect 88149 99451 88215 99454
rect 88517 99451 88583 99454
rect 97901 99451 97967 99454
rect 98678 99452 98684 99516
rect 98748 99514 98754 99516
rect 98821 99514 98887 99517
rect 98748 99512 98887 99514
rect 98748 99456 98826 99512
rect 98882 99456 98887 99512
rect 98748 99454 98887 99456
rect 101032 99514 101092 99893
rect 101446 99898 101632 99922
rect 101688 99898 101693 99954
rect 101811 99954 101877 99959
rect 101811 99924 101816 99954
rect 101872 99924 101877 99954
rect 101995 99954 102061 99959
rect 101446 99893 101693 99898
rect 101446 99862 101690 99893
rect 101446 99650 101506 99862
rect 101806 99860 101812 99924
rect 101876 99922 101882 99924
rect 101876 99862 101934 99922
rect 101995 99898 102000 99954
rect 102056 99922 102061 99954
rect 102547 99954 102613 99959
rect 102174 99922 102180 99924
rect 102056 99898 102180 99922
rect 101995 99893 102180 99898
rect 101998 99862 102180 99893
rect 101876 99860 101882 99862
rect 102174 99860 102180 99862
rect 102244 99860 102250 99924
rect 102547 99898 102552 99954
rect 102608 99898 102613 99954
rect 102547 99893 102613 99898
rect 102731 99954 102797 99959
rect 102731 99898 102736 99954
rect 102792 99898 102797 99954
rect 103099 99954 103165 99959
rect 102731 99893 102797 99898
rect 102550 99789 102610 99893
rect 102501 99784 102610 99789
rect 102501 99728 102506 99784
rect 102562 99728 102610 99784
rect 102501 99726 102610 99728
rect 102501 99723 102567 99726
rect 102734 99653 102794 99893
rect 102910 99860 102916 99924
rect 102980 99922 102986 99924
rect 103099 99922 103104 99954
rect 102980 99898 103104 99922
rect 103160 99898 103165 99954
rect 104939 99954 105005 99959
rect 103559 99922 103625 99925
rect 102980 99893 103165 99898
rect 103424 99920 103625 99922
rect 102980 99862 103162 99893
rect 103424 99864 103564 99920
rect 103620 99864 103625 99920
rect 104571 99920 104637 99925
rect 103424 99862 103625 99864
rect 102980 99860 102986 99862
rect 102869 99786 102935 99789
rect 103283 99788 103349 99789
rect 103278 99786 103284 99788
rect 102869 99784 102978 99786
rect 102869 99728 102874 99784
rect 102930 99728 102978 99784
rect 102869 99723 102978 99728
rect 103192 99726 103284 99786
rect 103278 99724 103284 99726
rect 103348 99724 103354 99788
rect 103424 99786 103484 99862
rect 103559 99859 103625 99862
rect 104203 99886 104269 99891
rect 104203 99830 104208 99886
rect 104264 99830 104269 99886
rect 104571 99864 104576 99920
rect 104632 99864 104637 99920
rect 104939 99898 104944 99954
rect 105000 99898 105005 99954
rect 106043 99954 106109 99959
rect 104939 99893 105005 99898
rect 104571 99859 104637 99864
rect 104203 99825 104269 99830
rect 103424 99726 103530 99786
rect 103283 99723 103349 99724
rect 101673 99650 101739 99653
rect 101446 99648 101739 99650
rect 101446 99592 101678 99648
rect 101734 99592 101739 99648
rect 101446 99590 101739 99592
rect 101673 99587 101739 99590
rect 101949 99648 102015 99653
rect 101949 99592 101954 99648
rect 102010 99592 102015 99648
rect 101949 99587 102015 99592
rect 102734 99648 102843 99653
rect 102734 99592 102782 99648
rect 102838 99592 102843 99648
rect 102734 99590 102843 99592
rect 102777 99587 102843 99590
rect 101397 99514 101463 99517
rect 101032 99512 101463 99514
rect 101032 99456 101402 99512
rect 101458 99456 101463 99512
rect 101032 99454 101463 99456
rect 98748 99452 98754 99454
rect 98821 99451 98887 99454
rect 101397 99451 101463 99454
rect 101622 99452 101628 99516
rect 101692 99514 101698 99516
rect 101952 99514 102012 99587
rect 101692 99454 102012 99514
rect 102317 99514 102383 99517
rect 102918 99514 102978 99723
rect 103470 99653 103530 99726
rect 104206 99653 104266 99825
rect 104574 99653 104634 99859
rect 104942 99789 105002 99893
rect 105302 99860 105308 99924
rect 105372 99922 105378 99924
rect 105583 99922 105649 99925
rect 106043 99924 106048 99954
rect 106104 99924 106109 99954
rect 107883 99954 107949 99959
rect 107377 99924 107443 99925
rect 105372 99920 105649 99922
rect 105372 99864 105588 99920
rect 105644 99864 105649 99920
rect 105372 99862 105649 99864
rect 105372 99860 105378 99862
rect 105583 99859 105649 99862
rect 106038 99860 106044 99924
rect 106108 99922 106114 99924
rect 107326 99922 107332 99924
rect 106108 99862 106166 99922
rect 107286 99862 107332 99922
rect 107396 99920 107443 99924
rect 107438 99864 107443 99920
rect 106108 99860 106114 99862
rect 107326 99860 107332 99862
rect 107396 99860 107443 99864
rect 107377 99859 107443 99860
rect 107515 99920 107581 99925
rect 107515 99864 107520 99920
rect 107576 99864 107581 99920
rect 107883 99898 107888 99954
rect 107944 99898 107949 99954
rect 108251 99954 108317 99959
rect 108251 99924 108256 99954
rect 108312 99924 108317 99954
rect 108619 99954 108728 99959
rect 107883 99893 107949 99898
rect 107515 99859 107581 99864
rect 107518 99789 107578 99859
rect 104942 99784 105051 99789
rect 104942 99728 104990 99784
rect 105046 99728 105051 99784
rect 104942 99726 105051 99728
rect 107518 99784 107627 99789
rect 107518 99728 107566 99784
rect 107622 99728 107627 99784
rect 107518 99726 107627 99728
rect 104985 99723 105051 99726
rect 107561 99723 107627 99726
rect 103094 99588 103100 99652
rect 103164 99650 103170 99652
rect 103329 99650 103395 99653
rect 103164 99648 103395 99650
rect 103164 99592 103334 99648
rect 103390 99592 103395 99648
rect 103164 99590 103395 99592
rect 103470 99648 103579 99653
rect 103470 99592 103518 99648
rect 103574 99592 103579 99648
rect 103470 99590 103579 99592
rect 103164 99588 103170 99590
rect 103329 99587 103395 99590
rect 103513 99587 103579 99590
rect 104157 99648 104266 99653
rect 104157 99592 104162 99648
rect 104218 99592 104266 99648
rect 104157 99590 104266 99592
rect 104525 99648 104634 99653
rect 104525 99592 104530 99648
rect 104586 99592 104634 99648
rect 104525 99590 104634 99592
rect 104801 99650 104867 99653
rect 107469 99652 107535 99653
rect 104801 99648 106474 99650
rect 104801 99592 104806 99648
rect 104862 99592 106474 99648
rect 104801 99590 106474 99592
rect 104157 99587 104223 99590
rect 104525 99587 104591 99590
rect 104801 99587 104867 99590
rect 102317 99512 102978 99514
rect 102317 99456 102322 99512
rect 102378 99456 102978 99512
rect 102317 99454 102978 99456
rect 106414 99514 106474 99590
rect 107469 99648 107516 99652
rect 107580 99650 107586 99652
rect 107469 99592 107474 99648
rect 107469 99588 107516 99592
rect 107580 99590 107626 99650
rect 107580 99588 107586 99590
rect 107469 99587 107535 99588
rect 107469 99514 107535 99517
rect 106414 99512 107535 99514
rect 106414 99456 107474 99512
rect 107530 99456 107535 99512
rect 106414 99454 107535 99456
rect 101692 99452 101698 99454
rect 102317 99451 102383 99454
rect 107469 99451 107535 99454
rect 107653 99514 107719 99517
rect 107886 99514 107946 99893
rect 108246 99860 108252 99924
rect 108316 99922 108322 99924
rect 108316 99862 108374 99922
rect 108619 99898 108624 99954
rect 108680 99898 108728 99954
rect 108619 99896 108728 99898
rect 108990 99922 109050 99998
rect 109174 99998 110644 100058
rect 109174 99922 109234 99998
rect 110638 99996 110644 99998
rect 110708 99996 110714 100060
rect 111750 100058 111810 100134
rect 115890 100134 124444 100194
rect 115890 100058 115950 100134
rect 124438 100132 124444 100134
rect 124508 100132 124514 100196
rect 111750 99998 115950 100058
rect 111379 99954 111445 99959
rect 108619 99893 108685 99896
rect 108803 99886 108869 99891
rect 108316 99860 108322 99862
rect 108803 99830 108808 99886
rect 108864 99830 108869 99886
rect 108990 99862 109234 99922
rect 109447 99922 109513 99925
rect 109447 99920 109786 99922
rect 109447 99864 109452 99920
rect 109508 99864 109786 99920
rect 109447 99862 109786 99864
rect 109447 99859 109513 99862
rect 108803 99825 108869 99830
rect 108062 99724 108068 99788
rect 108132 99786 108138 99788
rect 108389 99786 108455 99789
rect 108132 99784 108455 99786
rect 108132 99728 108394 99784
rect 108450 99728 108455 99784
rect 108132 99726 108455 99728
rect 108132 99724 108138 99726
rect 108389 99723 108455 99726
rect 108297 99652 108363 99653
rect 108246 99650 108252 99652
rect 108206 99590 108252 99650
rect 108316 99648 108363 99652
rect 108358 99592 108363 99648
rect 108246 99588 108252 99590
rect 108316 99588 108363 99592
rect 108430 99588 108436 99652
rect 108500 99650 108506 99652
rect 108665 99650 108731 99653
rect 108500 99648 108731 99650
rect 108500 99592 108670 99648
rect 108726 99592 108731 99648
rect 108500 99590 108731 99592
rect 108500 99588 108506 99590
rect 108297 99587 108363 99588
rect 108665 99587 108731 99590
rect 108806 99517 108866 99825
rect 107653 99512 107946 99514
rect 107653 99456 107658 99512
rect 107714 99456 107946 99512
rect 107653 99454 107946 99456
rect 108757 99512 108866 99517
rect 108757 99456 108762 99512
rect 108818 99456 108866 99512
rect 108757 99454 108866 99456
rect 109726 99514 109786 99862
rect 109902 99860 109908 99924
rect 109972 99922 109978 99924
rect 110183 99922 110249 99925
rect 109972 99920 110249 99922
rect 109972 99864 110188 99920
rect 110244 99864 110249 99920
rect 109972 99862 110249 99864
rect 109972 99860 109978 99862
rect 110183 99859 110249 99862
rect 111006 99860 111012 99924
rect 111076 99922 111082 99924
rect 111195 99922 111261 99925
rect 111076 99920 111261 99922
rect 111076 99864 111200 99920
rect 111256 99864 111261 99920
rect 111379 99898 111384 99954
rect 111440 99922 111445 99954
rect 116163 99954 116229 99959
rect 111558 99922 111564 99924
rect 111440 99898 111564 99922
rect 111379 99893 111564 99898
rect 111076 99862 111261 99864
rect 111382 99862 111564 99893
rect 111076 99860 111082 99862
rect 111195 99859 111261 99862
rect 111558 99860 111564 99862
rect 111628 99860 111634 99924
rect 111747 99920 111813 99925
rect 111747 99864 111752 99920
rect 111808 99864 111813 99920
rect 111747 99859 111813 99864
rect 113311 99922 113377 99925
rect 114507 99922 114573 99925
rect 113311 99920 113834 99922
rect 113311 99864 113316 99920
rect 113372 99864 113834 99920
rect 113311 99862 113834 99864
rect 113311 99859 113377 99862
rect 111750 99789 111810 99859
rect 110643 99784 110709 99789
rect 110643 99728 110648 99784
rect 110704 99728 110709 99784
rect 110643 99723 110709 99728
rect 111701 99784 111810 99789
rect 111701 99728 111706 99784
rect 111762 99728 111810 99784
rect 111701 99726 111810 99728
rect 111701 99723 111767 99726
rect 110646 99653 110706 99723
rect 110597 99648 110706 99653
rect 110597 99592 110602 99648
rect 110658 99592 110706 99648
rect 110597 99590 110706 99592
rect 112069 99650 112135 99653
rect 112069 99648 112178 99650
rect 112069 99592 112074 99648
rect 112130 99592 112178 99648
rect 110597 99587 110663 99590
rect 112069 99587 112178 99592
rect 111333 99514 111399 99517
rect 109726 99512 111399 99514
rect 109726 99456 111338 99512
rect 111394 99456 111399 99512
rect 109726 99454 111399 99456
rect 107653 99451 107719 99454
rect 108757 99451 108823 99454
rect 111333 99451 111399 99454
rect 83414 99388 83523 99393
rect 83414 99332 83462 99388
rect 83518 99332 83523 99388
rect 83414 99330 83523 99332
rect 83457 99327 83523 99330
rect 85062 99316 85068 99380
rect 85132 99378 85138 99380
rect 85205 99378 85271 99381
rect 85132 99376 85271 99378
rect 85132 99320 85210 99376
rect 85266 99320 85271 99376
rect 85132 99318 85271 99320
rect 85132 99316 85138 99318
rect 85205 99315 85271 99318
rect 111190 99316 111196 99380
rect 111260 99378 111266 99380
rect 111609 99378 111675 99381
rect 111260 99376 111675 99378
rect 111260 99320 111614 99376
rect 111670 99320 111675 99376
rect 111260 99318 111675 99320
rect 112118 99378 112178 99587
rect 113774 99514 113834 99862
rect 114507 99920 115306 99922
rect 114507 99864 114512 99920
rect 114568 99864 115306 99920
rect 116163 99898 116168 99954
rect 116224 99898 116229 99954
rect 116347 99954 116413 99959
rect 116347 99924 116352 99954
rect 116408 99924 116413 99954
rect 117083 99954 117149 99959
rect 116163 99893 116229 99898
rect 114507 99862 115306 99864
rect 114507 99859 114573 99862
rect 114134 99724 114140 99788
rect 114204 99786 114210 99788
rect 114323 99786 114389 99789
rect 114204 99784 114389 99786
rect 114204 99728 114328 99784
rect 114384 99728 114389 99784
rect 114204 99726 114389 99728
rect 114204 99724 114210 99726
rect 114323 99723 114389 99726
rect 114694 99750 115122 99786
rect 114694 99726 115018 99750
rect 114694 99653 114754 99726
rect 115013 99694 115018 99726
rect 115074 99694 115122 99750
rect 115013 99692 115122 99694
rect 115013 99689 115079 99692
rect 114645 99648 114754 99653
rect 114645 99592 114650 99648
rect 114706 99592 114754 99648
rect 114645 99590 114754 99592
rect 114645 99587 114711 99590
rect 113909 99514 113975 99517
rect 113774 99512 113975 99514
rect 113774 99456 113914 99512
rect 113970 99456 113975 99512
rect 113774 99454 113975 99456
rect 113909 99451 113975 99454
rect 115246 99393 115306 99862
rect 116166 99786 116226 99893
rect 116342 99860 116348 99924
rect 116412 99922 116418 99924
rect 116412 99862 116470 99922
rect 116531 99920 116597 99925
rect 117083 99924 117088 99954
rect 117144 99924 117149 99954
rect 118463 99954 118529 99959
rect 116531 99864 116536 99920
rect 116592 99864 116597 99920
rect 116412 99860 116418 99862
rect 116531 99859 116597 99864
rect 117078 99860 117084 99924
rect 117148 99922 117154 99924
rect 117148 99862 117206 99922
rect 117148 99860 117154 99862
rect 117814 99860 117820 99924
rect 117884 99922 117890 99924
rect 118279 99922 118345 99925
rect 117884 99920 118345 99922
rect 117884 99864 118284 99920
rect 118340 99864 118345 99920
rect 118463 99898 118468 99954
rect 118524 99898 118529 99954
rect 118463 99893 118529 99898
rect 118923 99954 118989 99959
rect 118923 99898 118928 99954
rect 118984 99898 118989 99954
rect 120395 99954 120461 99959
rect 118923 99893 118989 99898
rect 119751 99922 119817 99925
rect 119751 99920 120136 99922
rect 117884 99862 118345 99864
rect 117884 99860 117890 99862
rect 118279 99859 118345 99862
rect 116393 99786 116459 99789
rect 116166 99784 116459 99786
rect 116166 99728 116398 99784
rect 116454 99728 116459 99784
rect 116166 99726 116459 99728
rect 116393 99723 116459 99726
rect 116117 99514 116183 99517
rect 116534 99514 116594 99859
rect 118233 99788 118299 99789
rect 118182 99786 118188 99788
rect 118142 99726 118188 99786
rect 118252 99784 118299 99788
rect 118294 99728 118299 99784
rect 118182 99724 118188 99726
rect 118252 99724 118299 99728
rect 118233 99723 118299 99724
rect 116710 99588 116716 99652
rect 116780 99650 116786 99652
rect 117221 99650 117287 99653
rect 116780 99648 117287 99650
rect 116780 99592 117226 99648
rect 117282 99592 117287 99648
rect 116780 99590 117287 99592
rect 116780 99588 116786 99590
rect 117221 99587 117287 99590
rect 117998 99588 118004 99652
rect 118068 99650 118074 99652
rect 118466 99650 118526 99893
rect 118926 99786 118986 99893
rect 119751 99864 119756 99920
rect 119812 99864 120136 99920
rect 120395 99898 120400 99954
rect 120456 99898 120461 99954
rect 120763 99954 120829 99959
rect 121039 99956 121105 99959
rect 120763 99924 120768 99954
rect 120824 99924 120829 99954
rect 120996 99954 121105 99956
rect 120395 99893 120461 99898
rect 119751 99862 120136 99864
rect 119751 99859 119817 99862
rect 120076 99789 120136 99862
rect 118742 99726 118986 99786
rect 119613 99788 119679 99789
rect 119613 99784 119660 99788
rect 119724 99786 119730 99788
rect 119613 99728 119618 99784
rect 118742 99653 118802 99726
rect 119613 99724 119660 99728
rect 119724 99726 119770 99786
rect 120073 99784 120139 99789
rect 120073 99728 120078 99784
rect 120134 99728 120139 99784
rect 119724 99724 119730 99726
rect 119613 99723 119679 99724
rect 120073 99723 120139 99728
rect 118068 99590 118526 99650
rect 118693 99648 118802 99653
rect 118693 99592 118698 99648
rect 118754 99592 118802 99648
rect 118693 99590 118802 99592
rect 118068 99588 118074 99590
rect 118693 99587 118759 99590
rect 120398 99517 120458 99893
rect 120758 99860 120764 99924
rect 120828 99922 120834 99924
rect 120828 99862 120886 99922
rect 120996 99898 121044 99954
rect 121100 99898 121105 99954
rect 120996 99893 121105 99898
rect 121499 99954 121565 99959
rect 121499 99898 121504 99954
rect 121560 99898 121565 99954
rect 125639 99954 125705 99959
rect 121499 99893 121565 99898
rect 122051 99922 122117 99925
rect 122511 99922 122577 99925
rect 123891 99922 123957 99925
rect 124070 99922 124076 99924
rect 122051 99920 122252 99922
rect 120828 99860 120834 99862
rect 120996 99788 121056 99893
rect 120942 99724 120948 99788
rect 121012 99726 121056 99788
rect 121012 99724 121018 99726
rect 116117 99512 116594 99514
rect 116117 99456 116122 99512
rect 116178 99456 116594 99512
rect 116117 99454 116594 99456
rect 117221 99516 117287 99517
rect 117221 99512 117268 99516
rect 117332 99514 117338 99516
rect 117221 99456 117226 99512
rect 116117 99451 116183 99454
rect 117221 99452 117268 99456
rect 117332 99454 117378 99514
rect 120398 99512 120507 99517
rect 120398 99456 120446 99512
rect 120502 99456 120507 99512
rect 120398 99454 120507 99456
rect 121502 99514 121562 99893
rect 121683 99886 121749 99891
rect 121683 99830 121688 99886
rect 121744 99830 121749 99886
rect 122051 99864 122056 99920
rect 122112 99864 122252 99920
rect 122051 99862 122252 99864
rect 122051 99859 122117 99862
rect 121683 99825 121749 99830
rect 121686 99653 121746 99825
rect 122192 99653 122252 99862
rect 122511 99920 122620 99922
rect 122511 99864 122516 99920
rect 122572 99864 122620 99920
rect 122511 99859 122620 99864
rect 123891 99920 124076 99922
rect 123891 99864 123896 99920
rect 123952 99864 124076 99920
rect 123891 99862 124076 99864
rect 123891 99859 123957 99862
rect 124070 99860 124076 99862
rect 124140 99860 124146 99924
rect 124259 99920 124325 99925
rect 124259 99864 124264 99920
rect 124320 99864 124325 99920
rect 124259 99859 124325 99864
rect 124627 99920 124693 99925
rect 124627 99864 124632 99920
rect 124688 99864 124693 99920
rect 124627 99859 124693 99864
rect 124806 99860 124812 99924
rect 124876 99922 124882 99924
rect 125271 99922 125337 99925
rect 124876 99920 125337 99922
rect 124876 99864 125276 99920
rect 125332 99864 125337 99920
rect 125639 99898 125644 99954
rect 125700 99898 125705 99954
rect 125639 99893 125705 99898
rect 125915 99954 125981 99959
rect 126191 99956 126257 99959
rect 125915 99898 125920 99954
rect 125976 99898 125981 99954
rect 126148 99954 126257 99956
rect 126148 99924 126196 99954
rect 125915 99893 125981 99898
rect 124876 99862 125337 99864
rect 124876 99860 124882 99862
rect 125271 99859 125337 99862
rect 122419 99788 122485 99789
rect 122560 99788 122620 99859
rect 122414 99786 122420 99788
rect 122328 99726 122420 99786
rect 122414 99724 122420 99726
rect 122484 99724 122490 99788
rect 122560 99726 122604 99788
rect 122598 99724 122604 99726
rect 122668 99724 122674 99788
rect 122419 99723 122485 99724
rect 121637 99648 121746 99653
rect 121637 99592 121642 99648
rect 121698 99592 121746 99648
rect 121637 99590 121746 99592
rect 122189 99648 122255 99653
rect 122189 99592 122194 99648
rect 122250 99592 122255 99648
rect 121637 99587 121703 99590
rect 122189 99587 122255 99592
rect 124262 99650 124322 99859
rect 124397 99650 124463 99653
rect 124262 99648 124463 99650
rect 124262 99592 124402 99648
rect 124458 99592 124463 99648
rect 124262 99590 124463 99592
rect 124397 99587 124463 99590
rect 122097 99514 122163 99517
rect 121502 99512 122163 99514
rect 121502 99456 122102 99512
rect 122158 99456 122163 99512
rect 121502 99454 122163 99456
rect 124630 99514 124690 99859
rect 125501 99514 125567 99517
rect 124630 99512 125567 99514
rect 124630 99456 125506 99512
rect 125562 99456 125567 99512
rect 124630 99454 125567 99456
rect 125642 99514 125702 99893
rect 125918 99653 125978 99893
rect 126094 99860 126100 99924
rect 126164 99898 126196 99924
rect 126252 99898 126257 99954
rect 126164 99893 126257 99898
rect 126467 99954 126533 99959
rect 126467 99898 126472 99954
rect 126528 99898 126533 99954
rect 126651 99954 126717 99959
rect 126651 99924 126656 99954
rect 126712 99924 126717 99954
rect 126467 99893 126533 99898
rect 126164 99862 126208 99893
rect 126164 99860 126170 99862
rect 125869 99648 125978 99653
rect 126237 99650 126303 99653
rect 125869 99592 125874 99648
rect 125930 99592 125978 99648
rect 125869 99590 125978 99592
rect 126102 99648 126303 99650
rect 126102 99592 126242 99648
rect 126298 99592 126303 99648
rect 126102 99590 126303 99592
rect 125869 99587 125935 99590
rect 125777 99514 125843 99517
rect 125642 99512 125843 99514
rect 125642 99456 125782 99512
rect 125838 99456 125843 99512
rect 125642 99454 125843 99456
rect 117332 99452 117338 99454
rect 117221 99451 117287 99452
rect 120441 99451 120507 99454
rect 122097 99451 122163 99454
rect 125501 99451 125567 99454
rect 125777 99451 125843 99454
rect 115197 99388 115306 99393
rect 112253 99378 112319 99381
rect 112118 99376 112319 99378
rect 112118 99320 112258 99376
rect 112314 99320 112319 99376
rect 115197 99332 115202 99388
rect 115258 99332 115306 99388
rect 115197 99330 115306 99332
rect 125593 99378 125659 99381
rect 126102 99378 126162 99590
rect 126237 99587 126303 99590
rect 125593 99376 126162 99378
rect 115197 99327 115263 99330
rect 112118 99318 112319 99320
rect 111260 99316 111266 99318
rect 111609 99315 111675 99318
rect 112253 99315 112319 99318
rect 125593 99320 125598 99376
rect 125654 99320 126162 99376
rect 125593 99318 126162 99320
rect 125593 99315 125659 99318
rect 126145 99242 126211 99245
rect 126470 99242 126530 99893
rect 126646 99860 126652 99924
rect 126716 99922 126722 99924
rect 126716 99862 126774 99922
rect 126716 99860 126722 99862
rect 126145 99240 126530 99242
rect 126145 99184 126150 99240
rect 126206 99184 126530 99240
rect 126145 99182 126530 99184
rect 126145 99179 126211 99182
rect 89294 98364 89300 98428
rect 89364 98426 89370 98428
rect 89897 98426 89963 98429
rect 89364 98424 89963 98426
rect 89364 98368 89902 98424
rect 89958 98368 89963 98424
rect 89364 98366 89963 98368
rect 89364 98364 89370 98366
rect 89897 98363 89963 98366
rect 100150 98364 100156 98428
rect 100220 98426 100226 98428
rect 100661 98426 100727 98429
rect 100220 98424 100727 98426
rect 100220 98368 100666 98424
rect 100722 98368 100727 98424
rect 100220 98366 100727 98368
rect 100220 98364 100226 98366
rect 100661 98363 100727 98366
rect 122046 98364 122052 98428
rect 122116 98426 122122 98428
rect 122557 98426 122623 98429
rect 122116 98424 122623 98426
rect 122116 98368 122562 98424
rect 122618 98368 122623 98424
rect 122116 98366 122623 98368
rect 122116 98364 122122 98366
rect 122557 98363 122623 98366
rect 84193 98290 84259 98293
rect 84326 98290 84332 98292
rect 84193 98288 84332 98290
rect 84193 98232 84198 98288
rect 84254 98232 84332 98288
rect 84193 98230 84332 98232
rect 84193 98227 84259 98230
rect 84326 98228 84332 98230
rect 84396 98228 84402 98292
rect 85665 98290 85731 98293
rect 85798 98290 85804 98292
rect 85665 98288 85804 98290
rect 85665 98232 85670 98288
rect 85726 98232 85804 98288
rect 85665 98230 85804 98232
rect 85665 98227 85731 98230
rect 85798 98228 85804 98230
rect 85868 98228 85874 98292
rect 86350 98228 86356 98292
rect 86420 98290 86426 98292
rect 86493 98290 86559 98293
rect 86420 98288 86559 98290
rect 86420 98232 86498 98288
rect 86554 98232 86559 98288
rect 86420 98230 86559 98232
rect 86420 98228 86426 98230
rect 86493 98227 86559 98230
rect 90030 98228 90036 98292
rect 90100 98290 90106 98292
rect 90173 98290 90239 98293
rect 93393 98292 93459 98293
rect 93342 98290 93348 98292
rect 90100 98288 90239 98290
rect 90100 98232 90178 98288
rect 90234 98232 90239 98288
rect 90100 98230 90239 98232
rect 93302 98230 93348 98290
rect 93412 98288 93459 98292
rect 93454 98232 93459 98288
rect 90100 98228 90106 98230
rect 90173 98227 90239 98230
rect 93342 98228 93348 98230
rect 93412 98228 93459 98232
rect 95182 98228 95188 98292
rect 95252 98290 95258 98292
rect 95325 98290 95391 98293
rect 95252 98288 95391 98290
rect 95252 98232 95330 98288
rect 95386 98232 95391 98288
rect 95252 98230 95391 98232
rect 95252 98228 95258 98230
rect 93393 98227 93459 98228
rect 95325 98227 95391 98230
rect 99966 98228 99972 98292
rect 100036 98290 100042 98292
rect 100201 98290 100267 98293
rect 101765 98292 101831 98293
rect 101765 98290 101812 98292
rect 100036 98288 100267 98290
rect 100036 98232 100206 98288
rect 100262 98232 100267 98288
rect 100036 98230 100267 98232
rect 101720 98288 101812 98290
rect 101720 98232 101770 98288
rect 101720 98230 101812 98232
rect 100036 98228 100042 98230
rect 100201 98227 100267 98230
rect 101765 98228 101812 98230
rect 101876 98228 101882 98292
rect 102041 98290 102107 98293
rect 102174 98290 102180 98292
rect 102041 98288 102180 98290
rect 102041 98232 102046 98288
rect 102102 98232 102180 98288
rect 102041 98230 102180 98232
rect 101765 98227 101831 98228
rect 102041 98227 102107 98230
rect 102174 98228 102180 98230
rect 102244 98228 102250 98292
rect 102910 98228 102916 98292
rect 102980 98290 102986 98292
rect 103053 98290 103119 98293
rect 102980 98288 103119 98290
rect 102980 98232 103058 98288
rect 103114 98232 103119 98288
rect 102980 98230 103119 98232
rect 102980 98228 102986 98230
rect 103053 98227 103119 98230
rect 103605 98292 103671 98293
rect 105261 98292 105327 98293
rect 103605 98288 103652 98292
rect 103716 98290 103722 98292
rect 105261 98290 105308 98292
rect 103605 98232 103610 98288
rect 103605 98228 103652 98232
rect 103716 98230 103762 98290
rect 105216 98288 105308 98290
rect 105216 98232 105266 98288
rect 105216 98230 105308 98232
rect 103716 98228 103722 98230
rect 105261 98228 105308 98230
rect 105372 98228 105378 98292
rect 122782 98228 122788 98292
rect 122852 98290 122858 98292
rect 124029 98290 124095 98293
rect 126053 98292 126119 98293
rect 126053 98290 126100 98292
rect 122852 98288 124095 98290
rect 122852 98232 124034 98288
rect 124090 98232 124095 98288
rect 122852 98230 124095 98232
rect 126008 98288 126100 98290
rect 126008 98232 126058 98288
rect 126008 98230 126100 98232
rect 122852 98228 122858 98230
rect 103605 98227 103671 98228
rect 105261 98227 105327 98228
rect 124029 98227 124095 98230
rect 126053 98228 126100 98230
rect 126164 98228 126170 98292
rect 126462 98228 126468 98292
rect 126532 98290 126538 98292
rect 126881 98290 126947 98293
rect 126532 98288 126947 98290
rect 126532 98232 126886 98288
rect 126942 98232 126947 98288
rect 126532 98230 126947 98232
rect 126532 98228 126538 98230
rect 126053 98227 126119 98228
rect 126881 98227 126947 98230
rect 91318 98092 91324 98156
rect 91388 98154 91394 98156
rect 92197 98154 92263 98157
rect 91388 98152 92263 98154
rect 91388 98096 92202 98152
rect 92258 98096 92263 98152
rect 91388 98094 92263 98096
rect 91388 98092 91394 98094
rect 92197 98091 92263 98094
rect 100334 98092 100340 98156
rect 100404 98154 100410 98156
rect 100569 98154 100635 98157
rect 100404 98152 100635 98154
rect 100404 98096 100574 98152
rect 100630 98096 100635 98152
rect 100404 98094 100635 98096
rect 100404 98092 100410 98094
rect 100569 98091 100635 98094
rect 110086 98092 110092 98156
rect 110156 98154 110162 98156
rect 110321 98154 110387 98157
rect 126697 98156 126763 98157
rect 126646 98154 126652 98156
rect 110156 98152 110387 98154
rect 110156 98096 110326 98152
rect 110382 98096 110387 98152
rect 110156 98094 110387 98096
rect 126606 98094 126652 98154
rect 126716 98152 126763 98156
rect 126758 98096 126763 98152
rect 110156 98092 110162 98094
rect 110321 98091 110387 98094
rect 126646 98092 126652 98094
rect 126716 98092 126763 98096
rect 126697 98091 126763 98092
rect 89621 98018 89687 98021
rect 92289 98018 92355 98021
rect 89621 98016 92355 98018
rect 89621 97960 89626 98016
rect 89682 97960 92294 98016
rect 92350 97960 92355 98016
rect 89621 97958 92355 97960
rect 89621 97955 89687 97958
rect 92289 97955 92355 97958
rect 89110 97820 89116 97884
rect 89180 97882 89186 97884
rect 89621 97882 89687 97885
rect 89180 97880 89687 97882
rect 89180 97824 89626 97880
rect 89682 97824 89687 97880
rect 89180 97822 89687 97824
rect 89180 97820 89186 97822
rect 89621 97819 89687 97822
rect 94814 97820 94820 97884
rect 94884 97882 94890 97884
rect 95141 97882 95207 97885
rect 94884 97880 95207 97882
rect 94884 97824 95146 97880
rect 95202 97824 95207 97880
rect 94884 97822 95207 97824
rect 94884 97820 94890 97822
rect 95141 97819 95207 97822
rect 98637 97746 98703 97749
rect 122966 97746 122972 97748
rect 98637 97744 122972 97746
rect 98637 97688 98642 97744
rect 98698 97688 122972 97744
rect 98637 97686 122972 97688
rect 98637 97683 98703 97686
rect 122966 97684 122972 97686
rect 123036 97684 123042 97748
rect 83958 97548 83964 97612
rect 84028 97610 84034 97612
rect 93117 97610 93183 97613
rect 84028 97608 93183 97610
rect 84028 97552 93122 97608
rect 93178 97552 93183 97608
rect 84028 97550 93183 97552
rect 84028 97548 84034 97550
rect 93117 97547 93183 97550
rect 95734 97548 95740 97612
rect 95804 97610 95810 97612
rect 96521 97610 96587 97613
rect 95804 97608 96587 97610
rect 95804 97552 96526 97608
rect 96582 97552 96587 97608
rect 95804 97550 96587 97552
rect 95804 97548 95810 97550
rect 96521 97547 96587 97550
rect 97533 97612 97599 97613
rect 98177 97612 98243 97613
rect 98913 97612 98979 97613
rect 97533 97608 97580 97612
rect 97644 97610 97650 97612
rect 97533 97552 97538 97608
rect 97533 97548 97580 97552
rect 97644 97550 97690 97610
rect 97644 97548 97650 97550
rect 98126 97548 98132 97612
rect 98196 97610 98243 97612
rect 98862 97610 98868 97612
rect 98196 97608 98288 97610
rect 98238 97552 98288 97608
rect 98196 97550 98288 97552
rect 98822 97550 98868 97610
rect 98932 97608 98979 97612
rect 98974 97552 98979 97608
rect 98196 97548 98243 97550
rect 98862 97548 98868 97550
rect 98932 97548 98979 97552
rect 97533 97547 97599 97548
rect 98177 97547 98243 97548
rect 98913 97547 98979 97548
rect 99097 97610 99163 97613
rect 99230 97610 99236 97612
rect 99097 97608 99236 97610
rect 99097 97552 99102 97608
rect 99158 97552 99236 97608
rect 99097 97550 99236 97552
rect 99097 97547 99163 97550
rect 99230 97548 99236 97550
rect 99300 97548 99306 97612
rect 113909 97610 113975 97613
rect 113909 97608 114570 97610
rect 113909 97552 113914 97608
rect 113970 97552 114570 97608
rect 113909 97550 114570 97552
rect 113909 97547 113975 97550
rect 97390 97412 97396 97476
rect 97460 97474 97466 97476
rect 97625 97474 97691 97477
rect 97460 97472 97691 97474
rect 97460 97416 97630 97472
rect 97686 97416 97691 97472
rect 97460 97414 97691 97416
rect 97460 97412 97466 97414
rect 97625 97411 97691 97414
rect 99005 97476 99071 97477
rect 99005 97472 99052 97476
rect 99116 97474 99122 97476
rect 99005 97416 99010 97472
rect 99005 97412 99052 97416
rect 99116 97414 99162 97474
rect 99116 97412 99122 97414
rect 99005 97411 99071 97412
rect 97206 97140 97212 97204
rect 97276 97202 97282 97204
rect 97809 97202 97875 97205
rect 97276 97200 97875 97202
rect 97276 97144 97814 97200
rect 97870 97144 97875 97200
rect 97276 97142 97875 97144
rect 97276 97140 97282 97142
rect 97809 97139 97875 97142
rect 98085 97066 98151 97069
rect 99782 97066 99788 97068
rect 98085 97064 99788 97066
rect 98085 97008 98090 97064
rect 98146 97008 99788 97064
rect 98085 97006 99788 97008
rect 98085 97003 98151 97006
rect 99782 97004 99788 97006
rect 99852 97004 99858 97068
rect 112478 97004 112484 97068
rect 112548 97066 112554 97068
rect 112989 97066 113055 97069
rect 112548 97064 113055 97066
rect 112548 97008 112994 97064
rect 113050 97008 113055 97064
rect 112548 97006 113055 97008
rect 112548 97004 112554 97006
rect 112989 97003 113055 97006
rect 112805 96930 112871 96933
rect 113030 96930 113036 96932
rect 112805 96928 113036 96930
rect 112805 96872 112810 96928
rect 112866 96872 113036 96928
rect 112805 96870 113036 96872
rect 112805 96867 112871 96870
rect 113030 96868 113036 96870
rect 113100 96868 113106 96932
rect 113582 96868 113588 96932
rect 113652 96930 113658 96932
rect 114369 96930 114435 96933
rect 113652 96928 114435 96930
rect 113652 96872 114374 96928
rect 114430 96872 114435 96928
rect 113652 96870 114435 96872
rect 113652 96868 113658 96870
rect 114369 96867 114435 96870
rect 106733 96794 106799 96797
rect 106460 96792 106799 96794
rect 106460 96736 106738 96792
rect 106794 96736 106799 96792
rect 106460 96734 106799 96736
rect 106460 96661 106520 96734
rect 106733 96731 106799 96734
rect 109350 96732 109356 96796
rect 109420 96794 109426 96796
rect 110229 96794 110295 96797
rect 112713 96796 112779 96797
rect 112662 96794 112668 96796
rect 109420 96792 110295 96794
rect 109420 96736 110234 96792
rect 110290 96736 110295 96792
rect 109420 96734 110295 96736
rect 112622 96734 112668 96794
rect 112732 96792 112779 96796
rect 112774 96736 112779 96792
rect 109420 96732 109426 96734
rect 110229 96731 110295 96734
rect 112662 96732 112668 96734
rect 112732 96732 112779 96736
rect 113950 96732 113956 96796
rect 114020 96794 114026 96796
rect 114185 96794 114251 96797
rect 114020 96792 114251 96794
rect 114020 96736 114190 96792
rect 114246 96736 114251 96792
rect 114020 96734 114251 96736
rect 114020 96732 114026 96734
rect 112713 96731 112779 96732
rect 114185 96731 114251 96734
rect 114369 96794 114435 96797
rect 114510 96794 114570 97550
rect 122966 97548 122972 97612
rect 123036 97610 123042 97612
rect 123937 97610 124003 97613
rect 123036 97608 124003 97610
rect 123036 97552 123942 97608
rect 123998 97552 124003 97608
rect 123036 97550 124003 97552
rect 123036 97548 123042 97550
rect 123937 97547 124003 97550
rect 116761 97474 116827 97477
rect 116894 97474 116900 97476
rect 116761 97472 116900 97474
rect 116761 97416 116766 97472
rect 116822 97416 116900 97472
rect 116761 97414 116900 97416
rect 116761 97411 116827 97414
rect 116894 97412 116900 97414
rect 116964 97412 116970 97476
rect 120993 97338 121059 97341
rect 121126 97338 121132 97340
rect 120993 97336 121132 97338
rect 120993 97280 120998 97336
rect 121054 97280 121132 97336
rect 120993 97278 121132 97280
rect 120993 97275 121059 97278
rect 121126 97276 121132 97278
rect 121196 97276 121202 97340
rect 126605 97338 126671 97341
rect 126830 97338 126836 97340
rect 126605 97336 126836 97338
rect 126605 97280 126610 97336
rect 126666 97280 126836 97336
rect 126605 97278 126836 97280
rect 126605 97275 126671 97278
rect 126830 97276 126836 97278
rect 126900 97276 126906 97340
rect 118417 97202 118483 97205
rect 119797 97204 119863 97205
rect 118550 97202 118556 97204
rect 118417 97200 118556 97202
rect 118417 97144 118422 97200
rect 118478 97144 118556 97200
rect 118417 97142 118556 97144
rect 118417 97139 118483 97142
rect 118550 97140 118556 97142
rect 118620 97140 118626 97204
rect 119797 97200 119844 97204
rect 119908 97202 119914 97204
rect 119797 97144 119802 97200
rect 119797 97140 119844 97144
rect 119908 97142 119954 97202
rect 119908 97140 119914 97142
rect 120574 97140 120580 97204
rect 120644 97202 120650 97204
rect 121085 97202 121151 97205
rect 120644 97200 121151 97202
rect 120644 97144 121090 97200
rect 121146 97144 121151 97200
rect 120644 97142 121151 97144
rect 120644 97140 120650 97142
rect 119797 97139 119863 97140
rect 121085 97139 121151 97142
rect 118233 97066 118299 97069
rect 118366 97066 118372 97068
rect 118233 97064 118372 97066
rect 118233 97008 118238 97064
rect 118294 97008 118372 97064
rect 118233 97006 118372 97008
rect 118233 97003 118299 97006
rect 118366 97004 118372 97006
rect 118436 97004 118442 97068
rect 120758 97066 120764 97068
rect 120582 97006 120764 97066
rect 120582 96933 120642 97006
rect 120758 97004 120764 97006
rect 120828 97004 120834 97068
rect 124990 97004 124996 97068
rect 125060 97066 125066 97068
rect 125409 97066 125475 97069
rect 125060 97064 125475 97066
rect 125060 97008 125414 97064
rect 125470 97008 125475 97064
rect 125060 97006 125475 97008
rect 125060 97004 125066 97006
rect 125409 97003 125475 97006
rect 116342 96868 116348 96932
rect 116412 96930 116418 96932
rect 118325 96930 118391 96933
rect 116412 96928 118391 96930
rect 116412 96872 118330 96928
rect 118386 96872 118391 96928
rect 116412 96870 118391 96872
rect 120582 96928 120691 96933
rect 120582 96872 120630 96928
rect 120686 96872 120691 96928
rect 120582 96870 120691 96872
rect 116412 96868 116418 96870
rect 118325 96867 118391 96870
rect 120625 96867 120691 96870
rect 120758 96868 120764 96932
rect 120828 96930 120834 96932
rect 121177 96930 121243 96933
rect 120828 96928 121243 96930
rect 120828 96872 121182 96928
rect 121238 96872 121243 96928
rect 120828 96870 121243 96872
rect 120828 96868 120834 96870
rect 121177 96867 121243 96870
rect 115657 96796 115723 96797
rect 114369 96792 114570 96794
rect 114369 96736 114374 96792
rect 114430 96736 114570 96792
rect 114369 96734 114570 96736
rect 114369 96731 114435 96734
rect 115606 96732 115612 96796
rect 115676 96794 115723 96796
rect 115676 96792 115768 96794
rect 115718 96736 115768 96792
rect 115676 96734 115768 96736
rect 115676 96732 115723 96734
rect 122230 96732 122236 96796
rect 122300 96794 122306 96796
rect 122649 96794 122715 96797
rect 122300 96792 122715 96794
rect 122300 96736 122654 96792
rect 122710 96736 122715 96792
rect 122300 96734 122715 96736
rect 122300 96732 122306 96734
rect 115657 96731 115723 96732
rect 122649 96731 122715 96734
rect 125225 96794 125291 96797
rect 125358 96794 125364 96796
rect 125225 96792 125364 96794
rect 125225 96736 125230 96792
rect 125286 96736 125364 96792
rect 125225 96734 125364 96736
rect 125225 96731 125291 96734
rect 125358 96732 125364 96734
rect 125428 96732 125434 96796
rect 106457 96656 106523 96661
rect 106457 96600 106462 96656
rect 106518 96600 106523 96656
rect 106457 96595 106523 96600
rect 108757 96660 108823 96661
rect 112897 96660 112963 96661
rect 108757 96656 108804 96660
rect 108868 96658 108874 96660
rect 112846 96658 112852 96660
rect 108757 96600 108762 96656
rect 108757 96596 108804 96600
rect 108868 96598 108914 96658
rect 112806 96598 112852 96658
rect 112916 96656 112963 96660
rect 112958 96600 112963 96656
rect 108868 96596 108874 96598
rect 112846 96596 112852 96598
rect 112916 96596 112963 96600
rect 113766 96596 113772 96660
rect 113836 96658 113842 96660
rect 114001 96658 114067 96661
rect 113836 96656 114067 96658
rect 113836 96600 114006 96656
rect 114062 96600 114067 96656
rect 113836 96598 114067 96600
rect 113836 96596 113842 96598
rect 108757 96595 108823 96596
rect 112897 96595 112963 96596
rect 114001 96595 114067 96598
rect 115565 96658 115631 96661
rect 115790 96658 115796 96660
rect 115565 96656 115796 96658
rect 115565 96600 115570 96656
rect 115626 96600 115796 96656
rect 115565 96598 115796 96600
rect 115565 96595 115631 96598
rect 115790 96596 115796 96598
rect 115860 96596 115866 96660
rect 125174 96596 125180 96660
rect 125244 96658 125250 96660
rect 125317 96658 125383 96661
rect 125244 96656 125383 96658
rect 125244 96600 125322 96656
rect 125378 96600 125383 96656
rect 125244 96598 125383 96600
rect 125244 96596 125250 96598
rect 125317 96595 125383 96598
rect 104249 96524 104315 96525
rect 104198 96522 104204 96524
rect 104158 96462 104204 96522
rect 104268 96520 104315 96524
rect 104310 96464 104315 96520
rect 104198 96460 104204 96462
rect 104268 96460 104315 96464
rect 104249 96459 104315 96460
rect 110413 96522 110479 96525
rect 111006 96522 111012 96524
rect 110413 96520 111012 96522
rect 110413 96464 110418 96520
rect 110474 96464 111012 96520
rect 110413 96462 111012 96464
rect 110413 96459 110479 96462
rect 111006 96460 111012 96462
rect 111076 96460 111082 96524
rect 82486 96324 82492 96388
rect 82556 96386 82562 96388
rect 97533 96386 97599 96389
rect 82556 96384 97599 96386
rect 82556 96328 97538 96384
rect 97594 96328 97599 96384
rect 82556 96326 97599 96328
rect 82556 96324 82562 96326
rect 97533 96323 97599 96326
rect 107142 96324 107148 96388
rect 107212 96386 107218 96388
rect 107285 96386 107351 96389
rect 107212 96384 107351 96386
rect 107212 96328 107290 96384
rect 107346 96328 107351 96384
rect 107212 96326 107351 96328
rect 107212 96324 107218 96326
rect 107285 96323 107351 96326
rect 111006 96324 111012 96388
rect 111076 96386 111082 96388
rect 111701 96386 111767 96389
rect 111076 96384 111767 96386
rect 111076 96328 111706 96384
rect 111762 96328 111767 96384
rect 111076 96326 111767 96328
rect 111076 96324 111082 96326
rect 111701 96323 111767 96326
rect 105118 96188 105124 96252
rect 105188 96250 105194 96252
rect 106089 96250 106155 96253
rect 105188 96248 106155 96250
rect 105188 96192 106094 96248
rect 106150 96192 106155 96248
rect 105188 96190 106155 96192
rect 105188 96188 105194 96190
rect 106089 96187 106155 96190
rect 106958 96188 106964 96252
rect 107028 96250 107034 96252
rect 107561 96250 107627 96253
rect 108665 96252 108731 96253
rect 108614 96250 108620 96252
rect 107028 96248 107627 96250
rect 107028 96192 107566 96248
rect 107622 96192 107627 96248
rect 107028 96190 107627 96192
rect 108574 96190 108620 96250
rect 108684 96248 108731 96252
rect 108726 96192 108731 96248
rect 107028 96188 107034 96190
rect 107561 96187 107627 96190
rect 108614 96188 108620 96190
rect 108684 96188 108731 96192
rect 109534 96188 109540 96252
rect 109604 96250 109610 96252
rect 110045 96250 110111 96253
rect 109604 96248 110111 96250
rect 109604 96192 110050 96248
rect 110106 96192 110111 96248
rect 109604 96190 110111 96192
rect 109604 96188 109610 96190
rect 108665 96187 108731 96188
rect 110045 96187 110111 96190
rect 119889 96114 119955 96117
rect 471973 96114 472039 96117
rect 119889 96112 472039 96114
rect 119889 96056 119894 96112
rect 119950 96056 471978 96112
rect 472034 96056 472039 96112
rect 119889 96054 472039 96056
rect 119889 96051 119955 96054
rect 471973 96051 472039 96054
rect 121545 95978 121611 95981
rect 488533 95978 488599 95981
rect 121545 95976 488599 95978
rect 121545 95920 121550 95976
rect 121606 95920 488538 95976
rect 488594 95920 488599 95976
rect 121545 95918 488599 95920
rect 121545 95915 121611 95918
rect 488533 95915 488599 95918
rect 122782 95780 122788 95844
rect 122852 95842 122858 95844
rect 521653 95842 521719 95845
rect 122852 95840 521719 95842
rect 122852 95784 521658 95840
rect 521714 95784 521719 95840
rect 122852 95782 521719 95784
rect 122852 95780 122858 95782
rect 521653 95779 521719 95782
rect 101765 95706 101831 95709
rect 101990 95706 101996 95708
rect 101765 95704 101996 95706
rect 101765 95648 101770 95704
rect 101826 95648 101996 95704
rect 101765 95646 101996 95648
rect 101765 95643 101831 95646
rect 101990 95644 101996 95646
rect 102060 95644 102066 95708
rect 104433 95706 104499 95709
rect 104566 95706 104572 95708
rect 104433 95704 104572 95706
rect 104433 95648 104438 95704
rect 104494 95648 104572 95704
rect 104433 95646 104572 95648
rect 104433 95643 104499 95646
rect 104566 95644 104572 95646
rect 104636 95644 104642 95708
rect 101806 95508 101812 95572
rect 101876 95570 101882 95572
rect 102041 95570 102107 95573
rect 101876 95568 102107 95570
rect 101876 95512 102046 95568
rect 102102 95512 102107 95568
rect 101876 95510 102107 95512
rect 101876 95508 101882 95510
rect 102041 95507 102107 95510
rect 102910 95508 102916 95572
rect 102980 95570 102986 95572
rect 103053 95570 103119 95573
rect 102980 95568 103119 95570
rect 102980 95512 103058 95568
rect 103114 95512 103119 95568
rect 102980 95510 103119 95512
rect 102980 95508 102986 95510
rect 103053 95507 103119 95510
rect 103646 95508 103652 95572
rect 103716 95570 103722 95572
rect 104065 95570 104131 95573
rect 103716 95568 104131 95570
rect 103716 95512 104070 95568
rect 104126 95512 104131 95568
rect 103716 95510 104131 95512
rect 103716 95508 103722 95510
rect 104065 95507 104131 95510
rect 104382 95508 104388 95572
rect 104452 95570 104458 95572
rect 104617 95570 104683 95573
rect 111425 95572 111491 95573
rect 111374 95570 111380 95572
rect 104452 95568 104683 95570
rect 104452 95512 104622 95568
rect 104678 95512 104683 95568
rect 104452 95510 104683 95512
rect 111334 95510 111380 95570
rect 111444 95568 111491 95572
rect 111486 95512 111491 95568
rect 104452 95508 104458 95510
rect 104617 95507 104683 95510
rect 111374 95508 111380 95510
rect 111444 95508 111491 95512
rect 111425 95507 111491 95508
rect 107745 95434 107811 95437
rect 108062 95434 108068 95436
rect 107745 95432 108068 95434
rect 107745 95376 107750 95432
rect 107806 95376 108068 95432
rect 107745 95374 108068 95376
rect 107745 95371 107811 95374
rect 108062 95372 108068 95374
rect 108132 95372 108138 95436
rect 93710 94692 93716 94756
rect 93780 94754 93786 94756
rect 153193 94754 153259 94757
rect 93780 94752 153259 94754
rect 93780 94696 153198 94752
rect 153254 94696 153259 94752
rect 93780 94694 153259 94696
rect 93780 94692 93786 94694
rect 153193 94691 153259 94694
rect 100518 94556 100524 94620
rect 100588 94618 100594 94620
rect 235993 94618 236059 94621
rect 100588 94616 236059 94618
rect 100588 94560 235998 94616
rect 236054 94560 236059 94616
rect 100588 94558 236059 94560
rect 100588 94556 100594 94558
rect 235993 94555 236059 94558
rect 104709 94482 104775 94485
rect 289813 94482 289879 94485
rect 104709 94480 289879 94482
rect 104709 94424 104714 94480
rect 104770 94424 289818 94480
rect 289874 94424 289879 94480
rect 104709 94422 289879 94424
rect 104709 94419 104775 94422
rect 289813 94419 289879 94422
rect 110638 93468 110644 93532
rect 110708 93530 110714 93532
rect 335353 93530 335419 93533
rect 110708 93528 335419 93530
rect 110708 93472 335358 93528
rect 335414 93472 335419 93528
rect 110708 93470 335419 93472
rect 110708 93468 110714 93470
rect 335353 93467 335419 93470
rect 110137 93394 110203 93397
rect 356053 93394 356119 93397
rect 110137 93392 356119 93394
rect 110137 93336 110142 93392
rect 110198 93336 356058 93392
rect 356114 93336 356119 93392
rect 110137 93334 356119 93336
rect 110137 93331 110203 93334
rect 356053 93331 356119 93334
rect 111558 93196 111564 93260
rect 111628 93258 111634 93260
rect 368473 93258 368539 93261
rect 111628 93256 368539 93258
rect 111628 93200 368478 93256
rect 368534 93200 368539 93256
rect 111628 93198 368539 93200
rect 111628 93196 111634 93198
rect 368473 93195 368539 93198
rect 112478 93060 112484 93124
rect 112548 93122 112554 93124
rect 389173 93122 389239 93125
rect 112548 93120 389239 93122
rect 112548 93064 389178 93120
rect 389234 93064 389239 93120
rect 112548 93062 389239 93064
rect 112548 93060 112554 93062
rect 389173 93059 389239 93062
rect -960 92714 480 92804
rect 3877 92714 3943 92717
rect -960 92712 3943 92714
rect -960 92656 3882 92712
rect 3938 92656 3943 92712
rect -960 92654 3943 92656
rect -960 92564 480 92654
rect 3877 92651 3943 92654
rect 124254 92380 124260 92444
rect 124324 92442 124330 92444
rect 125041 92442 125107 92445
rect 124324 92440 125107 92442
rect 124324 92384 125046 92440
rect 125102 92384 125107 92440
rect 124324 92382 125107 92384
rect 124324 92380 124330 92382
rect 125041 92379 125107 92382
rect 102726 91700 102732 91764
rect 102796 91762 102802 91764
rect 103145 91762 103211 91765
rect 102796 91760 103211 91762
rect 102796 91704 103150 91760
rect 103206 91704 103211 91760
rect 102796 91702 103211 91704
rect 102796 91700 102802 91702
rect 103145 91699 103211 91702
rect 115606 90748 115612 90812
rect 115676 90810 115682 90812
rect 420913 90810 420979 90813
rect 115676 90808 420979 90810
rect 115676 90752 420918 90808
rect 420974 90752 420979 90808
rect 115676 90750 420979 90752
rect 115676 90748 115682 90750
rect 420913 90747 420979 90750
rect 117262 90612 117268 90676
rect 117332 90674 117338 90676
rect 436093 90674 436159 90677
rect 117332 90672 436159 90674
rect 117332 90616 436098 90672
rect 436154 90616 436159 90672
rect 117332 90614 436159 90616
rect 117332 90612 117338 90614
rect 436093 90611 436159 90614
rect 120574 90476 120580 90540
rect 120644 90538 120650 90540
rect 485773 90538 485839 90541
rect 120644 90536 485839 90538
rect 120644 90480 485778 90536
rect 485834 90480 485839 90536
rect 120644 90478 485839 90480
rect 120644 90476 120650 90478
rect 485773 90475 485839 90478
rect 122598 90340 122604 90404
rect 122668 90402 122674 90404
rect 502333 90402 502399 90405
rect 122668 90400 502399 90402
rect 122668 90344 502338 90400
rect 502394 90344 502399 90400
rect 122668 90342 502399 90344
rect 122668 90340 122674 90342
rect 502333 90339 502399 90342
rect 94446 88980 94452 89044
rect 94516 89042 94522 89044
rect 98637 89042 98703 89045
rect 94516 89040 98703 89042
rect 94516 88984 98642 89040
rect 98698 88984 98703 89040
rect 94516 88982 98703 88984
rect 94516 88980 94522 88982
rect 98637 88979 98703 88982
rect 89294 88164 89300 88228
rect 89364 88226 89370 88228
rect 94497 88226 94563 88229
rect 89364 88224 94563 88226
rect 89364 88168 94502 88224
rect 94558 88168 94563 88224
rect 89364 88166 94563 88168
rect 89364 88164 89370 88166
rect 94497 88163 94563 88166
rect 59353 87546 59419 87549
rect 85798 87546 85804 87548
rect 59353 87544 85804 87546
rect 59353 87488 59358 87544
rect 59414 87488 85804 87544
rect 59353 87486 85804 87488
rect 59353 87483 59419 87486
rect 85798 87484 85804 87486
rect 85868 87484 85874 87548
rect 90582 87484 90588 87548
rect 90652 87546 90658 87548
rect 104433 87546 104499 87549
rect 90652 87544 104499 87546
rect 90652 87488 104438 87544
rect 104494 87488 104499 87544
rect 90652 87486 104499 87488
rect 90652 87484 90658 87486
rect 104433 87483 104499 87486
rect 580533 86050 580599 86053
rect 583520 86050 584960 86140
rect 580533 86048 584960 86050
rect 580533 85992 580538 86048
rect 580594 85992 584960 86048
rect 580533 85990 584960 85992
rect 580533 85987 580599 85990
rect 583520 85900 584960 85990
rect 102726 84900 102732 84964
rect 102796 84962 102802 84964
rect 270493 84962 270559 84965
rect 102796 84960 270559 84962
rect 102796 84904 270498 84960
rect 270554 84904 270559 84960
rect 102796 84902 270559 84904
rect 102796 84900 102802 84902
rect 270493 84899 270559 84902
rect 106038 84764 106044 84828
rect 106108 84826 106114 84828
rect 304993 84826 305059 84829
rect 106108 84824 305059 84826
rect 106108 84768 304998 84824
rect 305054 84768 305059 84824
rect 106108 84766 305059 84768
rect 106108 84764 106114 84766
rect 304993 84763 305059 84766
rect 124806 79324 124812 79388
rect 124876 79386 124882 79388
rect 535453 79386 535519 79389
rect 124876 79384 535519 79386
rect 124876 79328 535458 79384
rect 535514 79328 535519 79384
rect 124876 79326 535519 79328
rect 124876 79324 124882 79326
rect 535453 79323 535519 79326
rect -960 75986 480 76076
rect 3785 75986 3851 75989
rect -960 75984 3851 75986
rect -960 75928 3790 75984
rect 3846 75928 3851 75984
rect -960 75926 3851 75928
rect -960 75836 480 75926
rect 3785 75923 3851 75926
rect 579613 70410 579679 70413
rect 583520 70410 584960 70500
rect 579613 70408 584960 70410
rect 579613 70352 579618 70408
rect 579674 70352 584960 70408
rect 579613 70350 584960 70352
rect 579613 70347 579679 70350
rect 583520 70260 584960 70350
rect -960 59258 480 59348
rect 3693 59258 3759 59261
rect -960 59256 3759 59258
rect -960 59200 3698 59256
rect 3754 59200 3759 59256
rect -960 59198 3759 59200
rect -960 59108 480 59198
rect 3693 59195 3759 59198
rect 580441 54770 580507 54773
rect 583520 54770 584960 54860
rect 580441 54768 584960 54770
rect 580441 54712 580446 54768
rect 580502 54712 584960 54768
rect 580441 54710 584960 54712
rect 580441 54707 580507 54710
rect 583520 54620 584960 54710
rect -960 42530 480 42620
rect 3601 42530 3667 42533
rect -960 42528 3667 42530
rect -960 42472 3606 42528
rect 3662 42472 3667 42528
rect -960 42470 3667 42472
rect -960 42380 480 42470
rect 3601 42467 3667 42470
rect 93342 42060 93348 42124
rect 93412 42122 93418 42124
rect 157333 42122 157399 42125
rect 93412 42120 157399 42122
rect 93412 42064 157338 42120
rect 157394 42064 157399 42120
rect 93412 42062 157399 42064
rect 93412 42060 93418 42062
rect 157333 42059 157399 42062
rect 91318 40836 91324 40900
rect 91388 40898 91394 40900
rect 140773 40898 140839 40901
rect 91388 40896 140839 40898
rect 91388 40840 140778 40896
rect 140834 40840 140839 40896
rect 91388 40838 140839 40840
rect 91388 40836 91394 40838
rect 140773 40835 140839 40838
rect 94630 40700 94636 40764
rect 94700 40762 94706 40764
rect 169845 40762 169911 40765
rect 94700 40760 169911 40762
rect 94700 40704 169850 40760
rect 169906 40704 169911 40760
rect 94700 40702 169911 40704
rect 94700 40700 94706 40702
rect 169845 40699 169911 40702
rect 95734 40564 95740 40628
rect 95804 40626 95810 40628
rect 190453 40626 190519 40629
rect 95804 40624 190519 40626
rect 95804 40568 190458 40624
rect 190514 40568 190519 40624
rect 95804 40566 190519 40568
rect 95804 40564 95810 40566
rect 190453 40563 190519 40566
rect 108430 39340 108436 39404
rect 108500 39402 108506 39404
rect 336733 39402 336799 39405
rect 108500 39400 336799 39402
rect 108500 39344 336738 39400
rect 336794 39344 336799 39400
rect 108500 39342 336799 39344
rect 108500 39340 108506 39342
rect 336733 39339 336799 39342
rect 126278 39204 126284 39268
rect 126348 39266 126354 39268
rect 552013 39266 552079 39269
rect 126348 39264 552079 39266
rect 126348 39208 552018 39264
rect 552074 39208 552079 39264
rect 126348 39206 552079 39208
rect 126348 39204 126354 39206
rect 552013 39203 552079 39206
rect 583520 39130 584960 39220
rect 583342 39070 584960 39130
rect 583342 38994 583402 39070
rect 583520 38994 584960 39070
rect 583342 38980 584960 38994
rect 583342 38934 583586 38980
rect 128854 38660 128860 38724
rect 128924 38722 128930 38724
rect 583526 38722 583586 38934
rect 128924 38662 583586 38722
rect 128924 38660 128930 38662
rect 97206 38252 97212 38316
rect 97276 38314 97282 38316
rect 207013 38314 207079 38317
rect 97276 38312 207079 38314
rect 97276 38256 207018 38312
rect 207074 38256 207079 38312
rect 97276 38254 207079 38256
rect 97276 38252 97282 38254
rect 207013 38251 207079 38254
rect 98678 38116 98684 38180
rect 98748 38178 98754 38180
rect 223573 38178 223639 38181
rect 98748 38176 223639 38178
rect 98748 38120 223578 38176
rect 223634 38120 223639 38176
rect 98748 38118 223639 38120
rect 98748 38116 98754 38118
rect 223573 38115 223639 38118
rect 116710 37980 116716 38044
rect 116780 38042 116786 38044
rect 438853 38042 438919 38045
rect 116780 38040 438919 38042
rect 116780 37984 438858 38040
rect 438914 37984 438919 38040
rect 116780 37982 438919 37984
rect 116780 37980 116786 37982
rect 438853 37979 438919 37982
rect 117814 37844 117820 37908
rect 117884 37906 117890 37908
rect 451273 37906 451339 37909
rect 117884 37904 451339 37906
rect 117884 37848 451278 37904
rect 451334 37848 451339 37904
rect 117884 37846 451339 37848
rect 117884 37844 117890 37846
rect 451273 37843 451339 37846
rect 95918 37164 95924 37228
rect 95988 37226 95994 37228
rect 186313 37226 186379 37229
rect 95988 37224 186379 37226
rect 95988 37168 186318 37224
rect 186374 37168 186379 37224
rect 95988 37166 186379 37168
rect 95988 37164 95994 37166
rect 186313 37163 186379 37166
rect 97390 37028 97396 37092
rect 97460 37090 97466 37092
rect 202873 37090 202939 37093
rect 97460 37088 202939 37090
rect 97460 37032 202878 37088
rect 202934 37032 202939 37088
rect 97460 37030 202939 37032
rect 97460 37028 97466 37030
rect 202873 37027 202939 37030
rect 111190 36892 111196 36956
rect 111260 36954 111266 36956
rect 372613 36954 372679 36957
rect 111260 36952 372679 36954
rect 111260 36896 372618 36952
rect 372674 36896 372679 36952
rect 111260 36894 372679 36896
rect 111260 36892 111266 36894
rect 372613 36891 372679 36894
rect 112662 36756 112668 36820
rect 112732 36818 112738 36820
rect 385033 36818 385099 36821
rect 112732 36816 385099 36818
rect 112732 36760 385038 36816
rect 385094 36760 385099 36816
rect 112732 36758 385099 36760
rect 112732 36756 112738 36758
rect 385033 36755 385099 36758
rect 124990 36620 124996 36684
rect 125060 36682 125066 36684
rect 538213 36682 538279 36685
rect 125060 36680 538279 36682
rect 125060 36624 538218 36680
rect 538274 36624 538279 36680
rect 125060 36622 538279 36624
rect 125060 36620 125066 36622
rect 538213 36619 538279 36622
rect 126462 36484 126468 36548
rect 126532 36546 126538 36548
rect 554773 36546 554839 36549
rect 126532 36544 554839 36546
rect 126532 36488 554778 36544
rect 554834 36488 554839 36544
rect 126532 36486 554839 36488
rect 126532 36484 126538 36486
rect 554773 36483 554839 36486
rect 94814 36348 94820 36412
rect 94884 36410 94890 36412
rect 173893 36410 173959 36413
rect 94884 36408 173959 36410
rect 94884 36352 173898 36408
rect 173954 36352 173959 36408
rect 94884 36350 173959 36352
rect 94884 36348 94890 36350
rect 173893 36347 173959 36350
rect 116894 35668 116900 35732
rect 116964 35730 116970 35732
rect 434805 35730 434871 35733
rect 116964 35728 434871 35730
rect 116964 35672 434810 35728
rect 434866 35672 434871 35728
rect 116964 35670 434871 35672
rect 116964 35668 116970 35670
rect 434805 35667 434871 35670
rect 117078 35532 117084 35596
rect 117148 35594 117154 35596
rect 437473 35594 437539 35597
rect 117148 35592 437539 35594
rect 117148 35536 437478 35592
rect 437534 35536 437539 35592
rect 117148 35534 437539 35536
rect 117148 35532 117154 35534
rect 437473 35531 437539 35534
rect 118182 35396 118188 35460
rect 118252 35458 118258 35460
rect 451365 35458 451431 35461
rect 118252 35456 451431 35458
rect 118252 35400 451370 35456
rect 451426 35400 451431 35456
rect 118252 35398 451431 35400
rect 118252 35396 118258 35398
rect 451365 35395 451431 35398
rect 117998 35260 118004 35324
rect 118068 35322 118074 35324
rect 454033 35322 454099 35325
rect 118068 35320 454099 35322
rect 118068 35264 454038 35320
rect 454094 35264 454099 35320
rect 118068 35262 454099 35264
rect 118068 35260 118074 35262
rect 454033 35259 454099 35262
rect 120942 35124 120948 35188
rect 121012 35186 121018 35188
rect 484393 35186 484459 35189
rect 121012 35184 484459 35186
rect 121012 35128 484398 35184
rect 484454 35128 484459 35184
rect 121012 35126 484459 35128
rect 121012 35124 121018 35126
rect 484393 35123 484459 35126
rect 113582 33764 113588 33828
rect 113652 33826 113658 33828
rect 405733 33826 405799 33829
rect 113652 33824 405799 33826
rect 113652 33768 405738 33824
rect 405794 33768 405799 33824
rect 113652 33766 405799 33768
rect 113652 33764 113658 33766
rect 405733 33763 405799 33766
rect 113766 32540 113772 32604
rect 113836 32602 113842 32604
rect 401685 32602 401751 32605
rect 113836 32600 401751 32602
rect 113836 32544 401690 32600
rect 401746 32544 401751 32600
rect 113836 32542 401751 32544
rect 113836 32540 113842 32542
rect 401685 32539 401751 32542
rect 119654 32404 119660 32468
rect 119724 32466 119730 32468
rect 467925 32466 467991 32469
rect 119724 32464 467991 32466
rect 119724 32408 467930 32464
rect 467986 32408 467991 32464
rect 119724 32406 467991 32408
rect 119724 32404 119730 32406
rect 467925 32403 467991 32406
rect 107142 31044 107148 31108
rect 107212 31106 107218 31108
rect 318793 31106 318859 31109
rect 107212 31104 318859 31106
rect 107212 31048 318798 31104
rect 318854 31048 318859 31104
rect 107212 31046 318859 31048
rect 107212 31044 107218 31046
rect 318793 31043 318859 31046
rect 106958 30908 106964 30972
rect 107028 30970 107034 30972
rect 322933 30970 322999 30973
rect 107028 30968 322999 30970
rect 107028 30912 322938 30968
rect 322994 30912 322999 30968
rect 107028 30910 322999 30912
rect 107028 30908 107034 30910
rect 322933 30907 322999 30910
rect 105118 29548 105124 29612
rect 105188 29610 105194 29612
rect 306373 29610 306439 29613
rect 105188 29608 306439 29610
rect 105188 29552 306378 29608
rect 306434 29552 306439 29608
rect 105188 29550 306439 29552
rect 105188 29548 105194 29550
rect 306373 29547 306439 29550
rect 93526 28460 93532 28524
rect 93596 28522 93602 28524
rect 153285 28522 153351 28525
rect 93596 28520 153351 28522
rect 93596 28464 153290 28520
rect 153346 28464 153351 28520
rect 93596 28462 153351 28464
rect 93596 28460 93602 28462
rect 153285 28459 153351 28462
rect 104566 28324 104572 28388
rect 104636 28386 104642 28388
rect 285765 28386 285831 28389
rect 104636 28384 285831 28386
rect 104636 28328 285770 28384
rect 285826 28328 285831 28384
rect 104636 28326 285831 28328
rect 104636 28324 104642 28326
rect 285765 28323 285831 28326
rect 104382 28188 104388 28252
rect 104452 28250 104458 28252
rect 285673 28250 285739 28253
rect 104452 28248 285739 28250
rect 104452 28192 285678 28248
rect 285734 28192 285739 28248
rect 104452 28190 285739 28192
rect 104452 28188 104458 28190
rect 285673 28187 285739 28190
rect 100150 27100 100156 27164
rect 100220 27162 100226 27164
rect 240133 27162 240199 27165
rect 100220 27160 240199 27162
rect 100220 27104 240138 27160
rect 240194 27104 240199 27160
rect 100220 27102 240199 27104
rect 100220 27100 100226 27102
rect 240133 27099 240199 27102
rect 102910 26964 102916 27028
rect 102980 27026 102986 27028
rect 269113 27026 269179 27029
rect 102980 27024 269179 27026
rect 102980 26968 269118 27024
rect 269174 26968 269179 27024
rect 102980 26966 269179 26968
rect 102980 26964 102986 26966
rect 269113 26963 269179 26966
rect 103094 26828 103100 26892
rect 103164 26890 103170 26892
rect 273253 26890 273319 26893
rect 103164 26888 273319 26890
rect 103164 26832 273258 26888
rect 273314 26832 273319 26888
rect 103164 26830 273319 26832
rect 103164 26828 103170 26830
rect 273253 26827 273319 26830
rect -960 25802 480 25892
rect 3509 25802 3575 25805
rect -960 25800 3575 25802
rect -960 25744 3514 25800
rect 3570 25744 3575 25800
rect -960 25742 3575 25744
rect -960 25652 480 25742
rect 3509 25739 3575 25742
rect 101622 25468 101628 25532
rect 101692 25530 101698 25532
rect 255313 25530 255379 25533
rect 101692 25528 255379 25530
rect 101692 25472 255318 25528
rect 255374 25472 255379 25528
rect 101692 25470 255379 25472
rect 101692 25468 101698 25470
rect 255313 25467 255379 25470
rect 98862 24380 98868 24444
rect 98932 24442 98938 24444
rect 219433 24442 219499 24445
rect 98932 24440 219499 24442
rect 98932 24384 219438 24440
rect 219494 24384 219499 24440
rect 98932 24382 219499 24384
rect 98932 24380 98938 24382
rect 219433 24379 219499 24382
rect 108614 24244 108620 24308
rect 108684 24306 108690 24308
rect 339493 24306 339559 24309
rect 108684 24304 339559 24306
rect 108684 24248 339498 24304
rect 339554 24248 339559 24304
rect 108684 24246 339559 24248
rect 108684 24244 108690 24246
rect 339493 24243 339559 24246
rect 109350 24108 109356 24172
rect 109420 24170 109426 24172
rect 351913 24170 351979 24173
rect 109420 24168 351979 24170
rect 109420 24112 351918 24168
rect 351974 24112 351979 24168
rect 109420 24110 351979 24112
rect 109420 24108 109426 24110
rect 351913 24107 351979 24110
rect 580349 23490 580415 23493
rect 583520 23490 584960 23580
rect 580349 23488 584960 23490
rect 580349 23432 580354 23488
rect 580410 23432 584960 23488
rect 580349 23430 584960 23432
rect 580349 23427 580415 23430
rect 583520 23340 584960 23430
rect 101806 22884 101812 22948
rect 101876 22946 101882 22948
rect 256693 22946 256759 22949
rect 101876 22944 256759 22946
rect 101876 22888 256698 22944
rect 256754 22888 256759 22944
rect 101876 22886 256759 22888
rect 101876 22884 101882 22886
rect 256693 22883 256759 22886
rect 125174 22748 125180 22812
rect 125244 22810 125250 22812
rect 536833 22810 536899 22813
rect 125244 22808 536899 22810
rect 125244 22752 536838 22808
rect 536894 22752 536899 22808
rect 125244 22750 536899 22752
rect 125244 22748 125250 22750
rect 536833 22747 536899 22750
rect 126646 22612 126652 22676
rect 126716 22674 126722 22676
rect 553393 22674 553459 22677
rect 126716 22672 553459 22674
rect 126716 22616 553398 22672
rect 553454 22616 553459 22672
rect 126716 22614 553459 22616
rect 126716 22612 126722 22614
rect 553393 22611 553459 22614
rect 99046 21388 99052 21452
rect 99116 21450 99122 21452
rect 219525 21450 219591 21453
rect 99116 21448 219591 21450
rect 99116 21392 219530 21448
rect 219586 21392 219591 21448
rect 99116 21390 219591 21392
rect 99116 21388 99122 21390
rect 219525 21387 219591 21390
rect 122966 21252 122972 21316
rect 123036 21314 123042 21316
rect 520273 21314 520339 21317
rect 123036 21312 520339 21314
rect 123036 21256 520278 21312
rect 520334 21256 520339 21312
rect 123036 21254 520339 21256
rect 123036 21252 123042 21254
rect 520273 21251 520339 21254
rect 94998 20028 95004 20092
rect 95068 20090 95074 20092
rect 172513 20090 172579 20093
rect 95068 20088 172579 20090
rect 95068 20032 172518 20088
rect 172574 20032 172579 20088
rect 95068 20030 172579 20032
rect 95068 20028 95074 20030
rect 172513 20027 172579 20030
rect 126830 19892 126836 19956
rect 126900 19954 126906 19956
rect 550725 19954 550791 19957
rect 126900 19952 550791 19954
rect 126900 19896 550730 19952
rect 550786 19896 550791 19952
rect 126900 19894 550791 19896
rect 126900 19892 126906 19894
rect 550725 19891 550791 19894
rect 91502 18940 91508 19004
rect 91572 19002 91578 19004
rect 139393 19002 139459 19005
rect 91572 19000 139459 19002
rect 91572 18944 139398 19000
rect 139454 18944 139459 19000
rect 91572 18942 139459 18944
rect 91572 18940 91578 18942
rect 139393 18939 139459 18942
rect 119838 18804 119844 18868
rect 119908 18866 119914 18868
rect 470593 18866 470659 18869
rect 119908 18864 470659 18866
rect 119908 18808 470598 18864
rect 470654 18808 470659 18864
rect 119908 18806 470659 18808
rect 119908 18804 119914 18806
rect 470593 18803 470659 18806
rect 122230 18668 122236 18732
rect 122300 18730 122306 18732
rect 505093 18730 505159 18733
rect 122300 18728 505159 18730
rect 122300 18672 505098 18728
rect 505154 18672 505159 18728
rect 122300 18670 505159 18672
rect 122300 18668 122306 18670
rect 505093 18667 505159 18670
rect 125358 18532 125364 18596
rect 125428 18594 125434 18596
rect 534073 18594 534139 18597
rect 125428 18592 534139 18594
rect 125428 18536 534078 18592
rect 534134 18536 534139 18592
rect 125428 18534 534139 18536
rect 125428 18532 125434 18534
rect 534073 18531 534139 18534
rect 118366 17444 118372 17508
rect 118436 17506 118442 17508
rect 449893 17506 449959 17509
rect 118436 17504 449959 17506
rect 118436 17448 449898 17504
rect 449954 17448 449959 17504
rect 118436 17446 449959 17448
rect 118436 17444 118442 17446
rect 449893 17443 449959 17446
rect 118550 17308 118556 17372
rect 118620 17370 118626 17372
rect 452653 17370 452719 17373
rect 118620 17368 452719 17370
rect 118620 17312 452658 17368
rect 452714 17312 452719 17368
rect 118620 17310 452719 17312
rect 118620 17308 118626 17310
rect 452653 17307 452719 17310
rect 122414 17172 122420 17236
rect 122484 17234 122490 17236
rect 501045 17234 501111 17237
rect 122484 17232 501111 17234
rect 122484 17176 501050 17232
rect 501106 17176 501111 17232
rect 122484 17174 501111 17176
rect 122484 17172 122490 17174
rect 501045 17171 501111 17174
rect 113950 16084 113956 16148
rect 114020 16146 114026 16148
rect 403985 16146 404051 16149
rect 114020 16144 404051 16146
rect 114020 16088 403990 16144
rect 404046 16088 404051 16144
rect 114020 16086 404051 16088
rect 114020 16084 114026 16086
rect 403985 16083 404051 16086
rect 114134 15948 114140 16012
rect 114204 16010 114210 16012
rect 405089 16010 405155 16013
rect 114204 16008 405155 16010
rect 114204 15952 405094 16008
rect 405150 15952 405155 16008
rect 114204 15950 405155 15952
rect 114204 15948 114210 15950
rect 405089 15947 405155 15950
rect 115790 15812 115796 15876
rect 115860 15874 115866 15876
rect 420545 15874 420611 15877
rect 115860 15872 420611 15874
rect 115860 15816 420550 15872
rect 420606 15816 420611 15872
rect 115860 15814 420611 15816
rect 115860 15812 115866 15814
rect 420545 15811 420611 15814
rect 111374 14860 111380 14924
rect 111444 14922 111450 14924
rect 370865 14922 370931 14925
rect 111444 14920 370931 14922
rect 111444 14864 370870 14920
rect 370926 14864 370931 14920
rect 111444 14862 370931 14864
rect 111444 14860 111450 14862
rect 370865 14859 370931 14862
rect 111006 14724 111012 14788
rect 111076 14786 111082 14788
rect 371969 14786 372035 14789
rect 111076 14784 372035 14786
rect 111076 14728 371974 14784
rect 372030 14728 372035 14784
rect 111076 14726 372035 14728
rect 111076 14724 111082 14726
rect 371969 14723 372035 14726
rect 113030 14588 113036 14652
rect 113100 14650 113106 14652
rect 387425 14650 387491 14653
rect 113100 14648 387491 14650
rect 113100 14592 387430 14648
rect 387486 14592 387491 14648
rect 113100 14590 387491 14592
rect 113100 14588 113106 14590
rect 387425 14587 387491 14590
rect 112846 14452 112852 14516
rect 112916 14514 112922 14516
rect 388529 14514 388595 14517
rect 112916 14512 388595 14514
rect 112916 14456 388534 14512
rect 388590 14456 388595 14512
rect 112916 14454 388595 14456
rect 112916 14452 112922 14454
rect 388529 14451 388595 14454
rect 107326 13228 107332 13292
rect 107396 13290 107402 13292
rect 322289 13290 322355 13293
rect 107396 13288 322355 13290
rect 107396 13232 322294 13288
rect 322350 13232 322355 13288
rect 107396 13230 322355 13232
rect 107396 13228 107402 13230
rect 322289 13227 322355 13230
rect 108798 13092 108804 13156
rect 108868 13154 108874 13156
rect 338849 13154 338915 13157
rect 108868 13152 338915 13154
rect 108868 13096 338854 13152
rect 338910 13096 338915 13152
rect 108868 13094 338915 13096
rect 108868 13092 108874 13094
rect 338849 13091 338915 13094
rect 109534 12956 109540 13020
rect 109604 13018 109610 13020
rect 354305 13018 354371 13021
rect 109604 13016 354371 13018
rect 109604 12960 354310 13016
rect 354366 12960 354371 13016
rect 109604 12958 354371 12960
rect 109604 12956 109610 12958
rect 354305 12955 354371 12958
rect 93158 11732 93164 11796
rect 93228 11794 93234 11796
rect 156689 11794 156755 11797
rect 93228 11792 156755 11794
rect 93228 11736 156694 11792
rect 156750 11736 156755 11792
rect 93228 11734 156755 11736
rect 93228 11732 93234 11734
rect 156689 11731 156755 11734
rect 107510 11596 107516 11660
rect 107580 11658 107586 11660
rect 321185 11658 321251 11661
rect 107580 11656 321251 11658
rect 107580 11600 321190 11656
rect 321246 11600 321251 11656
rect 107580 11598 321251 11600
rect 107580 11596 107586 11598
rect 321185 11595 321251 11598
rect 103278 10372 103284 10436
rect 103348 10434 103354 10436
rect 272609 10434 272675 10437
rect 103348 10432 272675 10434
rect 103348 10376 272614 10432
rect 272670 10376 272675 10432
rect 103348 10374 272675 10376
rect 103348 10372 103354 10374
rect 272609 10371 272675 10374
rect 104198 10236 104204 10300
rect 104268 10298 104274 10300
rect 289169 10298 289235 10301
rect 104268 10296 289235 10298
rect 104268 10240 289174 10296
rect 289230 10240 289235 10296
rect 104268 10238 289235 10240
rect 104268 10236 104274 10238
rect 289169 10235 289235 10238
rect 97758 9420 97764 9484
rect 97828 9482 97834 9484
rect 203057 9482 203123 9485
rect 97828 9480 203123 9482
rect 97828 9424 203062 9480
rect 203118 9424 203123 9480
rect 97828 9422 203123 9424
rect 97828 9420 97834 9422
rect 203057 9419 203123 9422
rect 97574 9284 97580 9348
rect 97644 9346 97650 9348
rect 206369 9346 206435 9349
rect 97644 9344 206435 9346
rect 97644 9288 206374 9344
rect 206430 9288 206435 9344
rect 97644 9286 206435 9288
rect 97644 9284 97650 9286
rect 206369 9283 206435 9286
rect -960 9074 480 9164
rect 99966 9148 99972 9212
rect 100036 9210 100042 9212
rect 236177 9210 236243 9213
rect 100036 9208 236243 9210
rect 100036 9152 236182 9208
rect 236238 9152 236243 9208
rect 100036 9150 236243 9152
rect 100036 9148 100042 9150
rect 236177 9147 236243 9150
rect 3417 9074 3483 9077
rect -960 9072 3483 9074
rect -960 9016 3422 9072
rect 3478 9016 3483 9072
rect -960 9014 3483 9016
rect -960 8924 480 9014
rect 3417 9011 3483 9014
rect 100334 9012 100340 9076
rect 100404 9074 100410 9076
rect 239489 9074 239555 9077
rect 100404 9072 239555 9074
rect 100404 9016 239494 9072
rect 239550 9016 239555 9072
rect 100404 9014 239555 9016
rect 100404 9012 100410 9014
rect 239489 9011 239555 9014
rect 101990 8876 101996 8940
rect 102060 8938 102066 8940
rect 254945 8938 255011 8941
rect 102060 8936 255011 8938
rect 102060 8880 254950 8936
rect 255006 8880 255011 8936
rect 102060 8878 255011 8880
rect 102060 8876 102066 8878
rect 254945 8875 255011 8878
rect 580257 7850 580323 7853
rect 583520 7850 584960 7940
rect 580257 7848 584960 7850
rect 580257 7792 580262 7848
rect 580318 7792 584960 7848
rect 580257 7790 584960 7792
rect 580257 7787 580323 7790
rect 583520 7700 584960 7790
rect 42977 7578 43043 7581
rect 84326 7578 84332 7580
rect 42977 7576 84332 7578
rect 42977 7520 42982 7576
rect 43038 7520 84332 7576
rect 42977 7518 84332 7520
rect 42977 7515 43043 7518
rect 84326 7516 84332 7518
rect 84396 7516 84402 7580
rect 96102 7516 96108 7580
rect 96172 7578 96178 7580
rect 189809 7578 189875 7581
rect 96172 7576 189875 7578
rect 96172 7520 189814 7576
rect 189870 7520 189875 7576
rect 96172 7518 189875 7520
rect 96172 7516 96178 7518
rect 189809 7515 189875 7518
rect 99230 6564 99236 6628
rect 99300 6626 99306 6628
rect 222929 6626 222995 6629
rect 99300 6624 222995 6626
rect 99300 6568 222934 6624
rect 222990 6568 222995 6624
rect 99300 6566 222995 6568
rect 99300 6564 99306 6566
rect 222929 6563 222995 6566
rect 121126 6428 121132 6492
rect 121196 6490 121202 6492
rect 484577 6490 484643 6493
rect 121196 6488 484643 6490
rect 121196 6432 484582 6488
rect 484638 6432 484643 6488
rect 121196 6430 484643 6432
rect 121196 6428 121202 6430
rect 484577 6427 484643 6430
rect 120758 6292 120764 6356
rect 120828 6354 120834 6356
rect 487889 6354 487955 6357
rect 120828 6352 487955 6354
rect 120828 6296 487894 6352
rect 487950 6296 487955 6352
rect 120828 6294 487955 6296
rect 120828 6292 120834 6294
rect 487889 6291 487955 6294
rect 122046 6156 122052 6220
rect 122116 6218 122122 6220
rect 504449 6218 504515 6221
rect 122116 6216 504515 6218
rect 122116 6160 504454 6216
rect 504510 6160 504515 6216
rect 122116 6158 504515 6160
rect 122116 6156 122122 6158
rect 504449 6155 504515 6158
rect 59537 4994 59603 4997
rect 85614 4994 85620 4996
rect 59537 4992 85620 4994
rect 59537 4936 59542 4992
rect 59598 4936 85620 4992
rect 59537 4934 85620 4936
rect 59537 4931 59603 4934
rect 85614 4932 85620 4934
rect 85684 4932 85690 4996
rect 46289 4858 46355 4861
rect 83958 4858 83964 4860
rect 46289 4856 83964 4858
rect 46289 4800 46294 4856
rect 46350 4800 83964 4856
rect 46289 4798 83964 4800
rect 46289 4795 46355 4798
rect 83958 4796 83964 4798
rect 84028 4796 84034 4860
rect 90766 4796 90772 4860
rect 90836 4858 90842 4860
rect 122465 4858 122531 4861
rect 90836 4856 122531 4858
rect 90836 4800 122470 4856
rect 122526 4800 122531 4856
rect 90836 4798 122531 4800
rect 90836 4796 90842 4798
rect 122465 4795 122531 4798
rect 124070 4796 124076 4860
rect 124140 4858 124146 4860
rect 519905 4858 519971 4861
rect 124140 4856 519971 4858
rect 124140 4800 519910 4856
rect 519966 4800 519971 4856
rect 124140 4798 519971 4800
rect 124140 4796 124146 4798
rect 519905 4795 519971 4798
rect 89478 3436 89484 3500
rect 89548 3498 89554 3500
rect 105905 3498 105971 3501
rect 89548 3496 105971 3498
rect 89548 3440 105910 3496
rect 105966 3440 105971 3496
rect 89548 3438 105971 3440
rect 89548 3436 89554 3438
rect 105905 3435 105971 3438
rect 90950 3300 90956 3364
rect 91020 3362 91026 3364
rect 124673 3362 124739 3365
rect 91020 3360 124739 3362
rect 91020 3304 124678 3360
rect 124734 3304 124739 3360
rect 91020 3302 124739 3304
rect 91020 3300 91026 3302
rect 124673 3299 124739 3302
<< via3 >>
rect 122604 152628 122668 152692
rect 124260 152220 124324 152284
rect 83780 151948 83844 152012
rect 124444 151948 124508 152012
rect 82492 151812 82556 151876
rect 128860 150452 128924 150516
rect 83964 149364 84028 149428
rect 99788 100132 99852 100196
rect 83780 99996 83844 100060
rect 84148 99860 84212 99924
rect 85068 99920 85132 99924
rect 85068 99864 85072 99920
rect 85072 99864 85128 99920
rect 85128 99864 85132 99920
rect 85068 99860 85132 99864
rect 86356 99920 86420 99924
rect 86356 99864 86360 99920
rect 86360 99864 86416 99920
rect 86416 99864 86420 99920
rect 85620 99724 85684 99788
rect 86356 99860 86420 99864
rect 89116 99898 89120 99924
rect 89120 99898 89176 99924
rect 89176 99898 89180 99924
rect 89116 99860 89180 99898
rect 90036 99920 90100 99924
rect 90036 99864 90040 99920
rect 90040 99864 90096 99920
rect 90096 99864 90100 99920
rect 90036 99860 90100 99864
rect 90956 99898 90960 99924
rect 90960 99898 91016 99924
rect 91016 99898 91020 99924
rect 90956 99860 91020 99898
rect 90772 99784 90836 99788
rect 90772 99728 90776 99784
rect 90776 99728 90832 99784
rect 90832 99728 90836 99784
rect 90772 99724 90836 99728
rect 89484 99588 89548 99652
rect 90588 99588 90652 99652
rect 91508 99588 91572 99652
rect 93348 99860 93412 99924
rect 94452 99860 94516 99924
rect 95188 99860 95252 99924
rect 95924 99860 95988 99924
rect 93716 99724 93780 99788
rect 94636 99784 94700 99788
rect 94636 99728 94686 99784
rect 94686 99728 94700 99784
rect 94636 99724 94700 99728
rect 95004 99784 95068 99788
rect 95004 99728 95008 99784
rect 95008 99728 95064 99784
rect 95064 99728 95068 99784
rect 95004 99724 95068 99728
rect 96108 99724 96172 99788
rect 93532 99588 93596 99652
rect 98132 99860 98196 99924
rect 97764 99724 97828 99788
rect 100524 99860 100588 99924
rect 99788 99724 99852 99788
rect 98684 99452 98748 99516
rect 101812 99898 101816 99924
rect 101816 99898 101872 99924
rect 101872 99898 101876 99924
rect 101812 99860 101876 99898
rect 102180 99860 102244 99924
rect 102916 99860 102980 99924
rect 103284 99784 103348 99788
rect 103284 99728 103288 99784
rect 103288 99728 103344 99784
rect 103344 99728 103348 99784
rect 103284 99724 103348 99728
rect 101628 99452 101692 99516
rect 105308 99860 105372 99924
rect 106044 99898 106048 99924
rect 106048 99898 106104 99924
rect 106104 99898 106108 99924
rect 106044 99860 106108 99898
rect 107332 99920 107396 99924
rect 107332 99864 107382 99920
rect 107382 99864 107396 99920
rect 107332 99860 107396 99864
rect 103100 99588 103164 99652
rect 107516 99648 107580 99652
rect 107516 99592 107530 99648
rect 107530 99592 107580 99648
rect 107516 99588 107580 99592
rect 108252 99898 108256 99924
rect 108256 99898 108312 99924
rect 108312 99898 108316 99924
rect 108252 99860 108316 99898
rect 110644 99996 110708 100060
rect 124444 100132 124508 100196
rect 108068 99724 108132 99788
rect 108252 99648 108316 99652
rect 108252 99592 108302 99648
rect 108302 99592 108316 99648
rect 108252 99588 108316 99592
rect 108436 99588 108500 99652
rect 109908 99860 109972 99924
rect 111012 99860 111076 99924
rect 111564 99860 111628 99924
rect 85068 99316 85132 99380
rect 111196 99316 111260 99380
rect 114140 99724 114204 99788
rect 116348 99898 116352 99924
rect 116352 99898 116408 99924
rect 116408 99898 116412 99924
rect 116348 99860 116412 99898
rect 117084 99898 117088 99924
rect 117088 99898 117144 99924
rect 117144 99898 117148 99924
rect 117084 99860 117148 99898
rect 117820 99860 117884 99924
rect 118188 99784 118252 99788
rect 118188 99728 118238 99784
rect 118238 99728 118252 99784
rect 118188 99724 118252 99728
rect 116716 99588 116780 99652
rect 118004 99588 118068 99652
rect 119660 99784 119724 99788
rect 119660 99728 119674 99784
rect 119674 99728 119724 99784
rect 119660 99724 119724 99728
rect 120764 99898 120768 99924
rect 120768 99898 120824 99924
rect 120824 99898 120828 99924
rect 120764 99860 120828 99898
rect 120948 99724 121012 99788
rect 117268 99512 117332 99516
rect 117268 99456 117282 99512
rect 117282 99456 117332 99512
rect 117268 99452 117332 99456
rect 124076 99860 124140 99924
rect 124812 99860 124876 99924
rect 122420 99784 122484 99788
rect 122420 99728 122424 99784
rect 122424 99728 122480 99784
rect 122480 99728 122484 99784
rect 122420 99724 122484 99728
rect 122604 99724 122668 99788
rect 126100 99860 126164 99924
rect 126652 99898 126656 99924
rect 126656 99898 126712 99924
rect 126712 99898 126716 99924
rect 126652 99860 126716 99898
rect 89300 98364 89364 98428
rect 100156 98364 100220 98428
rect 122052 98364 122116 98428
rect 84332 98228 84396 98292
rect 85804 98228 85868 98292
rect 86356 98228 86420 98292
rect 90036 98228 90100 98292
rect 93348 98288 93412 98292
rect 93348 98232 93398 98288
rect 93398 98232 93412 98288
rect 93348 98228 93412 98232
rect 95188 98228 95252 98292
rect 99972 98228 100036 98292
rect 101812 98288 101876 98292
rect 101812 98232 101826 98288
rect 101826 98232 101876 98288
rect 101812 98228 101876 98232
rect 102180 98228 102244 98292
rect 102916 98228 102980 98292
rect 103652 98288 103716 98292
rect 103652 98232 103666 98288
rect 103666 98232 103716 98288
rect 103652 98228 103716 98232
rect 105308 98288 105372 98292
rect 105308 98232 105322 98288
rect 105322 98232 105372 98288
rect 105308 98228 105372 98232
rect 122788 98228 122852 98292
rect 126100 98288 126164 98292
rect 126100 98232 126114 98288
rect 126114 98232 126164 98288
rect 126100 98228 126164 98232
rect 126468 98228 126532 98292
rect 91324 98092 91388 98156
rect 100340 98092 100404 98156
rect 110092 98092 110156 98156
rect 126652 98152 126716 98156
rect 126652 98096 126702 98152
rect 126702 98096 126716 98152
rect 126652 98092 126716 98096
rect 89116 97820 89180 97884
rect 94820 97820 94884 97884
rect 122972 97684 123036 97748
rect 83964 97548 84028 97612
rect 95740 97548 95804 97612
rect 97580 97608 97644 97612
rect 97580 97552 97594 97608
rect 97594 97552 97644 97608
rect 97580 97548 97644 97552
rect 98132 97608 98196 97612
rect 98132 97552 98182 97608
rect 98182 97552 98196 97608
rect 98132 97548 98196 97552
rect 98868 97608 98932 97612
rect 98868 97552 98918 97608
rect 98918 97552 98932 97608
rect 98868 97548 98932 97552
rect 99236 97548 99300 97612
rect 97396 97412 97460 97476
rect 99052 97472 99116 97476
rect 99052 97416 99066 97472
rect 99066 97416 99116 97472
rect 99052 97412 99116 97416
rect 97212 97140 97276 97204
rect 99788 97004 99852 97068
rect 112484 97004 112548 97068
rect 113036 96868 113100 96932
rect 113588 96868 113652 96932
rect 109356 96732 109420 96796
rect 112668 96792 112732 96796
rect 112668 96736 112718 96792
rect 112718 96736 112732 96792
rect 112668 96732 112732 96736
rect 113956 96732 114020 96796
rect 122972 97548 123036 97612
rect 116900 97412 116964 97476
rect 121132 97276 121196 97340
rect 126836 97276 126900 97340
rect 118556 97140 118620 97204
rect 119844 97200 119908 97204
rect 119844 97144 119858 97200
rect 119858 97144 119908 97200
rect 119844 97140 119908 97144
rect 120580 97140 120644 97204
rect 118372 97004 118436 97068
rect 120764 97004 120828 97068
rect 124996 97004 125060 97068
rect 116348 96868 116412 96932
rect 120764 96868 120828 96932
rect 115612 96792 115676 96796
rect 115612 96736 115662 96792
rect 115662 96736 115676 96792
rect 115612 96732 115676 96736
rect 122236 96732 122300 96796
rect 125364 96732 125428 96796
rect 108804 96656 108868 96660
rect 108804 96600 108818 96656
rect 108818 96600 108868 96656
rect 108804 96596 108868 96600
rect 112852 96656 112916 96660
rect 112852 96600 112902 96656
rect 112902 96600 112916 96656
rect 112852 96596 112916 96600
rect 113772 96596 113836 96660
rect 115796 96596 115860 96660
rect 125180 96596 125244 96660
rect 104204 96520 104268 96524
rect 104204 96464 104254 96520
rect 104254 96464 104268 96520
rect 104204 96460 104268 96464
rect 111012 96460 111076 96524
rect 82492 96324 82556 96388
rect 107148 96324 107212 96388
rect 111012 96324 111076 96388
rect 105124 96188 105188 96252
rect 106964 96188 107028 96252
rect 108620 96248 108684 96252
rect 108620 96192 108670 96248
rect 108670 96192 108684 96248
rect 108620 96188 108684 96192
rect 109540 96188 109604 96252
rect 122788 95780 122852 95844
rect 101996 95644 102060 95708
rect 104572 95644 104636 95708
rect 101812 95508 101876 95572
rect 102916 95508 102980 95572
rect 103652 95508 103716 95572
rect 104388 95508 104452 95572
rect 111380 95568 111444 95572
rect 111380 95512 111430 95568
rect 111430 95512 111444 95568
rect 111380 95508 111444 95512
rect 108068 95372 108132 95436
rect 93716 94692 93780 94756
rect 100524 94556 100588 94620
rect 110644 93468 110708 93532
rect 111564 93196 111628 93260
rect 112484 93060 112548 93124
rect 124260 92380 124324 92444
rect 102732 91700 102796 91764
rect 115612 90748 115676 90812
rect 117268 90612 117332 90676
rect 120580 90476 120644 90540
rect 122604 90340 122668 90404
rect 94452 88980 94516 89044
rect 89300 88164 89364 88228
rect 85804 87484 85868 87548
rect 90588 87484 90652 87548
rect 102732 84900 102796 84964
rect 106044 84764 106108 84828
rect 124812 79324 124876 79388
rect 93348 42060 93412 42124
rect 91324 40836 91388 40900
rect 94636 40700 94700 40764
rect 95740 40564 95804 40628
rect 108436 39340 108500 39404
rect 126284 39204 126348 39268
rect 128860 38660 128924 38724
rect 97212 38252 97276 38316
rect 98684 38116 98748 38180
rect 116716 37980 116780 38044
rect 117820 37844 117884 37908
rect 95924 37164 95988 37228
rect 97396 37028 97460 37092
rect 111196 36892 111260 36956
rect 112668 36756 112732 36820
rect 124996 36620 125060 36684
rect 126468 36484 126532 36548
rect 94820 36348 94884 36412
rect 116900 35668 116964 35732
rect 117084 35532 117148 35596
rect 118188 35396 118252 35460
rect 118004 35260 118068 35324
rect 120948 35124 121012 35188
rect 113588 33764 113652 33828
rect 113772 32540 113836 32604
rect 119660 32404 119724 32468
rect 107148 31044 107212 31108
rect 106964 30908 107028 30972
rect 105124 29548 105188 29612
rect 93532 28460 93596 28524
rect 104572 28324 104636 28388
rect 104388 28188 104452 28252
rect 100156 27100 100220 27164
rect 102916 26964 102980 27028
rect 103100 26828 103164 26892
rect 101628 25468 101692 25532
rect 98868 24380 98932 24444
rect 108620 24244 108684 24308
rect 109356 24108 109420 24172
rect 101812 22884 101876 22948
rect 125180 22748 125244 22812
rect 126652 22612 126716 22676
rect 99052 21388 99116 21452
rect 122972 21252 123036 21316
rect 95004 20028 95068 20092
rect 126836 19892 126900 19956
rect 91508 18940 91572 19004
rect 119844 18804 119908 18868
rect 122236 18668 122300 18732
rect 125364 18532 125428 18596
rect 118372 17444 118436 17508
rect 118556 17308 118620 17372
rect 122420 17172 122484 17236
rect 113956 16084 114020 16148
rect 114140 15948 114204 16012
rect 115796 15812 115860 15876
rect 111380 14860 111444 14924
rect 111012 14724 111076 14788
rect 113036 14588 113100 14652
rect 112852 14452 112916 14516
rect 107332 13228 107396 13292
rect 108804 13092 108868 13156
rect 109540 12956 109604 13020
rect 93164 11732 93228 11796
rect 107516 11596 107580 11660
rect 103284 10372 103348 10436
rect 104204 10236 104268 10300
rect 97764 9420 97828 9484
rect 97580 9284 97644 9348
rect 99972 9148 100036 9212
rect 100340 9012 100404 9076
rect 101996 8876 102060 8940
rect 84332 7516 84396 7580
rect 96108 7516 96172 7580
rect 99236 6564 99300 6628
rect 121132 6428 121196 6492
rect 120764 6292 120828 6356
rect 122052 6156 122116 6220
rect 85620 4932 85684 4996
rect 83964 4796 84028 4860
rect 90772 4796 90836 4860
rect 124076 4796 124140 4860
rect 89484 3436 89548 3500
rect 90956 3300 91020 3364
<< metal4 >>
rect -9036 711868 -8416 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 -8416 711868
rect -9036 711548 -8416 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 -8416 711548
rect -9036 682954 -8416 711312
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 -8416 682954
rect -9036 682634 -8416 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 -8416 682634
rect -9036 646954 -8416 682398
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 -8416 646954
rect -9036 646634 -8416 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 -8416 646634
rect -9036 610954 -8416 646398
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 -8416 610954
rect -9036 610634 -8416 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 -8416 610634
rect -9036 574954 -8416 610398
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 -8416 574954
rect -9036 574634 -8416 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 -8416 574634
rect -9036 538954 -8416 574398
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 -8416 538954
rect -9036 538634 -8416 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 -8416 538634
rect -9036 502954 -8416 538398
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 -8416 502954
rect -9036 502634 -8416 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 -8416 502634
rect -9036 466954 -8416 502398
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 -8416 466954
rect -9036 466634 -8416 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 -8416 466634
rect -9036 430954 -8416 466398
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 -8416 430954
rect -9036 430634 -8416 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 -8416 430634
rect -9036 394954 -8416 430398
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 -8416 394954
rect -9036 394634 -8416 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 -8416 394634
rect -9036 358954 -8416 394398
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 -8416 358954
rect -9036 358634 -8416 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 -8416 358634
rect -9036 322954 -8416 358398
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 -8416 322954
rect -9036 322634 -8416 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 -8416 322634
rect -9036 286954 -8416 322398
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 -8416 286954
rect -9036 286634 -8416 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 -8416 286634
rect -9036 250954 -8416 286398
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 -8416 250954
rect -9036 250634 -8416 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 -8416 250634
rect -9036 214954 -8416 250398
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 -8416 214954
rect -9036 214634 -8416 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 -8416 214634
rect -9036 178954 -8416 214398
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 -8416 178954
rect -9036 178634 -8416 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 -8416 178634
rect -9036 142954 -8416 178398
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 -8416 142954
rect -9036 142634 -8416 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 -8416 142634
rect -9036 106954 -8416 142398
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 -8416 106954
rect -9036 106634 -8416 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 -8416 106634
rect -9036 70954 -8416 106398
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 -8416 70954
rect -9036 70634 -8416 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 -8416 70634
rect -9036 34954 -8416 70398
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 -8416 34954
rect -9036 34634 -8416 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 -8416 34634
rect -9036 -7376 -8416 34398
rect -8076 710908 -7456 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 -7456 710908
rect -8076 710588 -7456 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 -7456 710588
rect -8076 678454 -7456 710352
rect -8076 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 -7456 678454
rect -8076 678134 -7456 678218
rect -8076 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 -7456 678134
rect -8076 642454 -7456 677898
rect -8076 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 -7456 642454
rect -8076 642134 -7456 642218
rect -8076 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 -7456 642134
rect -8076 606454 -7456 641898
rect -8076 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 -7456 606454
rect -8076 606134 -7456 606218
rect -8076 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 -7456 606134
rect -8076 570454 -7456 605898
rect -8076 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 -7456 570454
rect -8076 570134 -7456 570218
rect -8076 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 -7456 570134
rect -8076 534454 -7456 569898
rect -8076 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 -7456 534454
rect -8076 534134 -7456 534218
rect -8076 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 -7456 534134
rect -8076 498454 -7456 533898
rect -8076 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 -7456 498454
rect -8076 498134 -7456 498218
rect -8076 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 -7456 498134
rect -8076 462454 -7456 497898
rect -8076 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 -7456 462454
rect -8076 462134 -7456 462218
rect -8076 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 -7456 462134
rect -8076 426454 -7456 461898
rect -8076 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 -7456 426454
rect -8076 426134 -7456 426218
rect -8076 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 -7456 426134
rect -8076 390454 -7456 425898
rect -8076 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 -7456 390454
rect -8076 390134 -7456 390218
rect -8076 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 -7456 390134
rect -8076 354454 -7456 389898
rect -8076 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 -7456 354454
rect -8076 354134 -7456 354218
rect -8076 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 -7456 354134
rect -8076 318454 -7456 353898
rect -8076 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 -7456 318454
rect -8076 318134 -7456 318218
rect -8076 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 -7456 318134
rect -8076 282454 -7456 317898
rect -8076 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 -7456 282454
rect -8076 282134 -7456 282218
rect -8076 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 -7456 282134
rect -8076 246454 -7456 281898
rect -8076 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 -7456 246454
rect -8076 246134 -7456 246218
rect -8076 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 -7456 246134
rect -8076 210454 -7456 245898
rect -8076 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 -7456 210454
rect -8076 210134 -7456 210218
rect -8076 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 -7456 210134
rect -8076 174454 -7456 209898
rect -8076 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 -7456 174454
rect -8076 174134 -7456 174218
rect -8076 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 -7456 174134
rect -8076 138454 -7456 173898
rect -8076 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 -7456 138454
rect -8076 138134 -7456 138218
rect -8076 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 -7456 138134
rect -8076 102454 -7456 137898
rect -8076 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 -7456 102454
rect -8076 102134 -7456 102218
rect -8076 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 -7456 102134
rect -8076 66454 -7456 101898
rect -8076 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 -7456 66454
rect -8076 66134 -7456 66218
rect -8076 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 -7456 66134
rect -8076 30454 -7456 65898
rect -8076 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 -7456 30454
rect -8076 30134 -7456 30218
rect -8076 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 -7456 30134
rect -8076 -6416 -7456 29898
rect -7116 709948 -6496 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 -6496 709948
rect -7116 709628 -6496 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 -6496 709628
rect -7116 673954 -6496 709392
rect -7116 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 -6496 673954
rect -7116 673634 -6496 673718
rect -7116 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 -6496 673634
rect -7116 637954 -6496 673398
rect -7116 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 -6496 637954
rect -7116 637634 -6496 637718
rect -7116 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 -6496 637634
rect -7116 601954 -6496 637398
rect -7116 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 -6496 601954
rect -7116 601634 -6496 601718
rect -7116 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 -6496 601634
rect -7116 565954 -6496 601398
rect -7116 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 -6496 565954
rect -7116 565634 -6496 565718
rect -7116 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 -6496 565634
rect -7116 529954 -6496 565398
rect -7116 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 -6496 529954
rect -7116 529634 -6496 529718
rect -7116 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 -6496 529634
rect -7116 493954 -6496 529398
rect -7116 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 -6496 493954
rect -7116 493634 -6496 493718
rect -7116 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 -6496 493634
rect -7116 457954 -6496 493398
rect -7116 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 -6496 457954
rect -7116 457634 -6496 457718
rect -7116 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 -6496 457634
rect -7116 421954 -6496 457398
rect -7116 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 -6496 421954
rect -7116 421634 -6496 421718
rect -7116 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 -6496 421634
rect -7116 385954 -6496 421398
rect -7116 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 -6496 385954
rect -7116 385634 -6496 385718
rect -7116 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 -6496 385634
rect -7116 349954 -6496 385398
rect -7116 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 -6496 349954
rect -7116 349634 -6496 349718
rect -7116 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 -6496 349634
rect -7116 313954 -6496 349398
rect -7116 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 -6496 313954
rect -7116 313634 -6496 313718
rect -7116 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 -6496 313634
rect -7116 277954 -6496 313398
rect -7116 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 -6496 277954
rect -7116 277634 -6496 277718
rect -7116 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 -6496 277634
rect -7116 241954 -6496 277398
rect -7116 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 -6496 241954
rect -7116 241634 -6496 241718
rect -7116 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 -6496 241634
rect -7116 205954 -6496 241398
rect -7116 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 -6496 205954
rect -7116 205634 -6496 205718
rect -7116 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 -6496 205634
rect -7116 169954 -6496 205398
rect -7116 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 -6496 169954
rect -7116 169634 -6496 169718
rect -7116 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 -6496 169634
rect -7116 133954 -6496 169398
rect -7116 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 -6496 133954
rect -7116 133634 -6496 133718
rect -7116 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 -6496 133634
rect -7116 97954 -6496 133398
rect -7116 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 -6496 97954
rect -7116 97634 -6496 97718
rect -7116 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 -6496 97634
rect -7116 61954 -6496 97398
rect -7116 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 -6496 61954
rect -7116 61634 -6496 61718
rect -7116 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 -6496 61634
rect -7116 25954 -6496 61398
rect -7116 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 -6496 25954
rect -7116 25634 -6496 25718
rect -7116 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 -6496 25634
rect -7116 -5456 -6496 25398
rect -6156 708988 -5536 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 -5536 708988
rect -6156 708668 -5536 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 -5536 708668
rect -6156 669454 -5536 708432
rect -6156 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 -5536 669454
rect -6156 669134 -5536 669218
rect -6156 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 -5536 669134
rect -6156 633454 -5536 668898
rect -6156 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 -5536 633454
rect -6156 633134 -5536 633218
rect -6156 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 -5536 633134
rect -6156 597454 -5536 632898
rect -6156 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 -5536 597454
rect -6156 597134 -5536 597218
rect -6156 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 -5536 597134
rect -6156 561454 -5536 596898
rect -6156 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 -5536 561454
rect -6156 561134 -5536 561218
rect -6156 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 -5536 561134
rect -6156 525454 -5536 560898
rect -6156 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 -5536 525454
rect -6156 525134 -5536 525218
rect -6156 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 -5536 525134
rect -6156 489454 -5536 524898
rect -6156 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 -5536 489454
rect -6156 489134 -5536 489218
rect -6156 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 -5536 489134
rect -6156 453454 -5536 488898
rect -6156 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 -5536 453454
rect -6156 453134 -5536 453218
rect -6156 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 -5536 453134
rect -6156 417454 -5536 452898
rect -6156 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 -5536 417454
rect -6156 417134 -5536 417218
rect -6156 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 -5536 417134
rect -6156 381454 -5536 416898
rect -6156 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 -5536 381454
rect -6156 381134 -5536 381218
rect -6156 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 -5536 381134
rect -6156 345454 -5536 380898
rect -6156 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 -5536 345454
rect -6156 345134 -5536 345218
rect -6156 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 -5536 345134
rect -6156 309454 -5536 344898
rect -6156 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 -5536 309454
rect -6156 309134 -5536 309218
rect -6156 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 -5536 309134
rect -6156 273454 -5536 308898
rect -6156 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 -5536 273454
rect -6156 273134 -5536 273218
rect -6156 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 -5536 273134
rect -6156 237454 -5536 272898
rect -6156 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 -5536 237454
rect -6156 237134 -5536 237218
rect -6156 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 -5536 237134
rect -6156 201454 -5536 236898
rect -6156 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 -5536 201454
rect -6156 201134 -5536 201218
rect -6156 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 -5536 201134
rect -6156 165454 -5536 200898
rect -6156 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 -5536 165454
rect -6156 165134 -5536 165218
rect -6156 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 -5536 165134
rect -6156 129454 -5536 164898
rect -6156 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 -5536 129454
rect -6156 129134 -5536 129218
rect -6156 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 -5536 129134
rect -6156 93454 -5536 128898
rect -6156 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 -5536 93454
rect -6156 93134 -5536 93218
rect -6156 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 -5536 93134
rect -6156 57454 -5536 92898
rect -6156 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 -5536 57454
rect -6156 57134 -5536 57218
rect -6156 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 -5536 57134
rect -6156 21454 -5536 56898
rect -6156 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 -5536 21454
rect -6156 21134 -5536 21218
rect -6156 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 -5536 21134
rect -6156 -4496 -5536 20898
rect -5196 708028 -4576 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 -4576 708028
rect -5196 707708 -4576 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 -4576 707708
rect -5196 700954 -4576 707472
rect -5196 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 -4576 700954
rect -5196 700634 -4576 700718
rect -5196 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 -4576 700634
rect -5196 664954 -4576 700398
rect -5196 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 -4576 664954
rect -5196 664634 -4576 664718
rect -5196 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 -4576 664634
rect -5196 628954 -4576 664398
rect -5196 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 -4576 628954
rect -5196 628634 -4576 628718
rect -5196 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 -4576 628634
rect -5196 592954 -4576 628398
rect -5196 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 -4576 592954
rect -5196 592634 -4576 592718
rect -5196 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 -4576 592634
rect -5196 556954 -4576 592398
rect -5196 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 -4576 556954
rect -5196 556634 -4576 556718
rect -5196 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 -4576 556634
rect -5196 520954 -4576 556398
rect -5196 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 -4576 520954
rect -5196 520634 -4576 520718
rect -5196 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 -4576 520634
rect -5196 484954 -4576 520398
rect -5196 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 -4576 484954
rect -5196 484634 -4576 484718
rect -5196 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 -4576 484634
rect -5196 448954 -4576 484398
rect -5196 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 -4576 448954
rect -5196 448634 -4576 448718
rect -5196 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 -4576 448634
rect -5196 412954 -4576 448398
rect -5196 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 -4576 412954
rect -5196 412634 -4576 412718
rect -5196 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 -4576 412634
rect -5196 376954 -4576 412398
rect -5196 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 -4576 376954
rect -5196 376634 -4576 376718
rect -5196 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 -4576 376634
rect -5196 340954 -4576 376398
rect -5196 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 -4576 340954
rect -5196 340634 -4576 340718
rect -5196 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 -4576 340634
rect -5196 304954 -4576 340398
rect -5196 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 -4576 304954
rect -5196 304634 -4576 304718
rect -5196 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 -4576 304634
rect -5196 268954 -4576 304398
rect -5196 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 -4576 268954
rect -5196 268634 -4576 268718
rect -5196 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 -4576 268634
rect -5196 232954 -4576 268398
rect -5196 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 -4576 232954
rect -5196 232634 -4576 232718
rect -5196 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 -4576 232634
rect -5196 196954 -4576 232398
rect -5196 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 -4576 196954
rect -5196 196634 -4576 196718
rect -5196 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 -4576 196634
rect -5196 160954 -4576 196398
rect -5196 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 -4576 160954
rect -5196 160634 -4576 160718
rect -5196 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 -4576 160634
rect -5196 124954 -4576 160398
rect -5196 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 -4576 124954
rect -5196 124634 -4576 124718
rect -5196 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 -4576 124634
rect -5196 88954 -4576 124398
rect -5196 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 -4576 88954
rect -5196 88634 -4576 88718
rect -5196 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 -4576 88634
rect -5196 52954 -4576 88398
rect -5196 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 -4576 52954
rect -5196 52634 -4576 52718
rect -5196 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 -4576 52634
rect -5196 16954 -4576 52398
rect -5196 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 -4576 16954
rect -5196 16634 -4576 16718
rect -5196 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 -4576 16634
rect -5196 -3536 -4576 16398
rect -4236 707068 -3616 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 -3616 707068
rect -4236 706748 -3616 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 -3616 706748
rect -4236 696454 -3616 706512
rect -4236 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 -3616 696454
rect -4236 696134 -3616 696218
rect -4236 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 -3616 696134
rect -4236 660454 -3616 695898
rect -4236 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 -3616 660454
rect -4236 660134 -3616 660218
rect -4236 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 -3616 660134
rect -4236 624454 -3616 659898
rect -4236 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 -3616 624454
rect -4236 624134 -3616 624218
rect -4236 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 -3616 624134
rect -4236 588454 -3616 623898
rect -4236 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 -3616 588454
rect -4236 588134 -3616 588218
rect -4236 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 -3616 588134
rect -4236 552454 -3616 587898
rect -4236 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 -3616 552454
rect -4236 552134 -3616 552218
rect -4236 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 -3616 552134
rect -4236 516454 -3616 551898
rect -4236 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 -3616 516454
rect -4236 516134 -3616 516218
rect -4236 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 -3616 516134
rect -4236 480454 -3616 515898
rect -4236 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 -3616 480454
rect -4236 480134 -3616 480218
rect -4236 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 -3616 480134
rect -4236 444454 -3616 479898
rect -4236 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 -3616 444454
rect -4236 444134 -3616 444218
rect -4236 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 -3616 444134
rect -4236 408454 -3616 443898
rect -4236 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 -3616 408454
rect -4236 408134 -3616 408218
rect -4236 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 -3616 408134
rect -4236 372454 -3616 407898
rect -4236 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 -3616 372454
rect -4236 372134 -3616 372218
rect -4236 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 -3616 372134
rect -4236 336454 -3616 371898
rect -4236 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 -3616 336454
rect -4236 336134 -3616 336218
rect -4236 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 -3616 336134
rect -4236 300454 -3616 335898
rect -4236 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 -3616 300454
rect -4236 300134 -3616 300218
rect -4236 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 -3616 300134
rect -4236 264454 -3616 299898
rect -4236 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 -3616 264454
rect -4236 264134 -3616 264218
rect -4236 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 -3616 264134
rect -4236 228454 -3616 263898
rect -4236 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 -3616 228454
rect -4236 228134 -3616 228218
rect -4236 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 -3616 228134
rect -4236 192454 -3616 227898
rect -4236 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 -3616 192454
rect -4236 192134 -3616 192218
rect -4236 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 -3616 192134
rect -4236 156454 -3616 191898
rect -4236 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 -3616 156454
rect -4236 156134 -3616 156218
rect -4236 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 -3616 156134
rect -4236 120454 -3616 155898
rect -4236 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 -3616 120454
rect -4236 120134 -3616 120218
rect -4236 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 -3616 120134
rect -4236 84454 -3616 119898
rect -4236 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 -3616 84454
rect -4236 84134 -3616 84218
rect -4236 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 -3616 84134
rect -4236 48454 -3616 83898
rect -4236 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 -3616 48454
rect -4236 48134 -3616 48218
rect -4236 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 -3616 48134
rect -4236 12454 -3616 47898
rect -4236 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 -3616 12454
rect -4236 12134 -3616 12218
rect -4236 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 -3616 12134
rect -4236 -2576 -3616 11898
rect -3276 706108 -2656 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 -2656 706108
rect -3276 705788 -2656 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 -2656 705788
rect -3276 691954 -2656 705552
rect -3276 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 -2656 691954
rect -3276 691634 -2656 691718
rect -3276 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 -2656 691634
rect -3276 655954 -2656 691398
rect -3276 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 -2656 655954
rect -3276 655634 -2656 655718
rect -3276 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 -2656 655634
rect -3276 619954 -2656 655398
rect -3276 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 -2656 619954
rect -3276 619634 -2656 619718
rect -3276 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 -2656 619634
rect -3276 583954 -2656 619398
rect -3276 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 -2656 583954
rect -3276 583634 -2656 583718
rect -3276 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 -2656 583634
rect -3276 547954 -2656 583398
rect -3276 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 -2656 547954
rect -3276 547634 -2656 547718
rect -3276 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 -2656 547634
rect -3276 511954 -2656 547398
rect -3276 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 -2656 511954
rect -3276 511634 -2656 511718
rect -3276 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 -2656 511634
rect -3276 475954 -2656 511398
rect -3276 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 -2656 475954
rect -3276 475634 -2656 475718
rect -3276 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 -2656 475634
rect -3276 439954 -2656 475398
rect -3276 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 -2656 439954
rect -3276 439634 -2656 439718
rect -3276 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 -2656 439634
rect -3276 403954 -2656 439398
rect -3276 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 -2656 403954
rect -3276 403634 -2656 403718
rect -3276 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 -2656 403634
rect -3276 367954 -2656 403398
rect -3276 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 -2656 367954
rect -3276 367634 -2656 367718
rect -3276 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 -2656 367634
rect -3276 331954 -2656 367398
rect -3276 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 -2656 331954
rect -3276 331634 -2656 331718
rect -3276 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 -2656 331634
rect -3276 295954 -2656 331398
rect -3276 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 -2656 295954
rect -3276 295634 -2656 295718
rect -3276 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 -2656 295634
rect -3276 259954 -2656 295398
rect -3276 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 -2656 259954
rect -3276 259634 -2656 259718
rect -3276 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 -2656 259634
rect -3276 223954 -2656 259398
rect -3276 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 -2656 223954
rect -3276 223634 -2656 223718
rect -3276 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 -2656 223634
rect -3276 187954 -2656 223398
rect -3276 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 -2656 187954
rect -3276 187634 -2656 187718
rect -3276 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 -2656 187634
rect -3276 151954 -2656 187398
rect -3276 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 -2656 151954
rect -3276 151634 -2656 151718
rect -3276 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 -2656 151634
rect -3276 115954 -2656 151398
rect -3276 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 -2656 115954
rect -3276 115634 -2656 115718
rect -3276 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 -2656 115634
rect -3276 79954 -2656 115398
rect -3276 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 -2656 79954
rect -3276 79634 -2656 79718
rect -3276 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 -2656 79634
rect -3276 43954 -2656 79398
rect -3276 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 -2656 43954
rect -3276 43634 -2656 43718
rect -3276 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 -2656 43634
rect -3276 7954 -2656 43398
rect -3276 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 -2656 7954
rect -3276 7634 -2656 7718
rect -3276 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 -2656 7634
rect -3276 -1616 -2656 7398
rect -2316 705148 -1696 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 -1696 705148
rect -2316 704828 -1696 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 -1696 704828
rect -2316 687454 -1696 704592
rect -2316 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 -1696 687454
rect -2316 687134 -1696 687218
rect -2316 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 -1696 687134
rect -2316 651454 -1696 686898
rect -2316 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 -1696 651454
rect -2316 651134 -1696 651218
rect -2316 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 -1696 651134
rect -2316 615454 -1696 650898
rect -2316 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 -1696 615454
rect -2316 615134 -1696 615218
rect -2316 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 -1696 615134
rect -2316 579454 -1696 614898
rect -2316 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 -1696 579454
rect -2316 579134 -1696 579218
rect -2316 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 -1696 579134
rect -2316 543454 -1696 578898
rect -2316 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 -1696 543454
rect -2316 543134 -1696 543218
rect -2316 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 -1696 543134
rect -2316 507454 -1696 542898
rect -2316 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 -1696 507454
rect -2316 507134 -1696 507218
rect -2316 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 -1696 507134
rect -2316 471454 -1696 506898
rect -2316 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 -1696 471454
rect -2316 471134 -1696 471218
rect -2316 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 -1696 471134
rect -2316 435454 -1696 470898
rect -2316 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 -1696 435454
rect -2316 435134 -1696 435218
rect -2316 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 -1696 435134
rect -2316 399454 -1696 434898
rect -2316 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 -1696 399454
rect -2316 399134 -1696 399218
rect -2316 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 -1696 399134
rect -2316 363454 -1696 398898
rect -2316 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 -1696 363454
rect -2316 363134 -1696 363218
rect -2316 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 -1696 363134
rect -2316 327454 -1696 362898
rect -2316 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 -1696 327454
rect -2316 327134 -1696 327218
rect -2316 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 -1696 327134
rect -2316 291454 -1696 326898
rect -2316 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 -1696 291454
rect -2316 291134 -1696 291218
rect -2316 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 -1696 291134
rect -2316 255454 -1696 290898
rect -2316 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 -1696 255454
rect -2316 255134 -1696 255218
rect -2316 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 -1696 255134
rect -2316 219454 -1696 254898
rect -2316 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 -1696 219454
rect -2316 219134 -1696 219218
rect -2316 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 -1696 219134
rect -2316 183454 -1696 218898
rect -2316 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 -1696 183454
rect -2316 183134 -1696 183218
rect -2316 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 -1696 183134
rect -2316 147454 -1696 182898
rect -2316 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 -1696 147454
rect -2316 147134 -1696 147218
rect -2316 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 -1696 147134
rect -2316 111454 -1696 146898
rect -2316 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 -1696 111454
rect -2316 111134 -1696 111218
rect -2316 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 -1696 111134
rect -2316 75454 -1696 110898
rect -2316 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 -1696 75454
rect -2316 75134 -1696 75218
rect -2316 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 -1696 75134
rect -2316 39454 -1696 74898
rect -2316 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 -1696 39454
rect -2316 39134 -1696 39218
rect -2316 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 -1696 39134
rect -2316 3454 -1696 38898
rect -2316 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 -1696 3454
rect -2316 3134 -1696 3218
rect -2316 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 -1696 3134
rect -2316 -656 -1696 2898
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 -1696 -656
rect -2316 -976 -1696 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 -1696 -976
rect -2316 -1244 -1696 -1212
rect 1794 705148 2414 711900
rect 1794 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 2414 705148
rect 1794 704828 2414 704912
rect 1794 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 2414 704828
rect 1794 687454 2414 704592
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -656 2414 2898
rect 1794 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 2414 -656
rect 1794 -976 2414 -892
rect 1794 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 2414 -976
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 -2656 -1616
rect -3276 -1936 -2656 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 -2656 -1936
rect -3276 -2204 -2656 -2172
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 -3616 -2576
rect -4236 -2896 -3616 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 -3616 -2896
rect -4236 -3164 -3616 -3132
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 -4576 -3536
rect -5196 -3856 -4576 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 -4576 -3856
rect -5196 -4124 -4576 -4092
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 -5536 -4496
rect -6156 -4816 -5536 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 -5536 -4816
rect -6156 -5084 -5536 -5052
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 -6496 -5456
rect -7116 -5776 -6496 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 -6496 -5776
rect -7116 -6044 -6496 -6012
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 -7456 -6416
rect -8076 -6736 -7456 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 -7456 -6736
rect -8076 -7004 -7456 -6972
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 -8416 -7376
rect -9036 -7696 -8416 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 -8416 -7696
rect -9036 -7964 -8416 -7932
rect 1794 -7964 2414 -1212
rect 6294 706108 6914 711900
rect 6294 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 6914 706108
rect 6294 705788 6914 705872
rect 6294 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 6914 705788
rect 6294 691954 6914 705552
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1616 6914 7398
rect 6294 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 6914 -1616
rect 6294 -1936 6914 -1852
rect 6294 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 6914 -1936
rect 6294 -7964 6914 -2172
rect 10794 707068 11414 711900
rect 10794 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 11414 707068
rect 10794 706748 11414 706832
rect 10794 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 11414 706748
rect 10794 696454 11414 706512
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2576 11414 11898
rect 10794 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 11414 -2576
rect 10794 -2896 11414 -2812
rect 10794 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 11414 -2896
rect 10794 -7964 11414 -3132
rect 15294 708028 15914 711900
rect 15294 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 15914 708028
rect 15294 707708 15914 707792
rect 15294 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 15914 707708
rect 15294 700954 15914 707472
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3536 15914 16398
rect 15294 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 15914 -3536
rect 15294 -3856 15914 -3772
rect 15294 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 15914 -3856
rect 15294 -7964 15914 -4092
rect 19794 708988 20414 711900
rect 19794 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 20414 708988
rect 19794 708668 20414 708752
rect 19794 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 20414 708668
rect 19794 669454 20414 708432
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4496 20414 20898
rect 19794 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 20414 -4496
rect 19794 -4816 20414 -4732
rect 19794 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 20414 -4816
rect 19794 -7964 20414 -5052
rect 24294 709948 24914 711900
rect 24294 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 24914 709948
rect 24294 709628 24914 709712
rect 24294 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 24914 709628
rect 24294 673954 24914 709392
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5456 24914 25398
rect 24294 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 24914 -5456
rect 24294 -5776 24914 -5692
rect 24294 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 24914 -5776
rect 24294 -7964 24914 -6012
rect 28794 710908 29414 711900
rect 28794 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 29414 710908
rect 28794 710588 29414 710672
rect 28794 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 29414 710588
rect 28794 678454 29414 710352
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6416 29414 29898
rect 28794 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 29414 -6416
rect 28794 -6736 29414 -6652
rect 28794 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 29414 -6736
rect 28794 -7964 29414 -6972
rect 33294 711868 33914 711900
rect 33294 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 33914 711868
rect 33294 711548 33914 711632
rect 33294 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 33914 711548
rect 33294 682954 33914 711312
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7376 33914 34398
rect 33294 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 33914 -7376
rect 33294 -7696 33914 -7612
rect 33294 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 33914 -7696
rect 33294 -7964 33914 -7932
rect 37794 705148 38414 711900
rect 37794 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 38414 705148
rect 37794 704828 38414 704912
rect 37794 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 38414 704828
rect 37794 687454 38414 704592
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -656 38414 2898
rect 37794 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 38414 -656
rect 37794 -976 38414 -892
rect 37794 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 38414 -976
rect 37794 -7964 38414 -1212
rect 42294 706108 42914 711900
rect 42294 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 42914 706108
rect 42294 705788 42914 705872
rect 42294 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 42914 705788
rect 42294 691954 42914 705552
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1616 42914 7398
rect 42294 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 42914 -1616
rect 42294 -1936 42914 -1852
rect 42294 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 42914 -1936
rect 42294 -7964 42914 -2172
rect 46794 707068 47414 711900
rect 46794 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 47414 707068
rect 46794 706748 47414 706832
rect 46794 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 47414 706748
rect 46794 696454 47414 706512
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2576 47414 11898
rect 46794 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 47414 -2576
rect 46794 -2896 47414 -2812
rect 46794 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 47414 -2896
rect 46794 -7964 47414 -3132
rect 51294 708028 51914 711900
rect 51294 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 51914 708028
rect 51294 707708 51914 707792
rect 51294 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 51914 707708
rect 51294 700954 51914 707472
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3536 51914 16398
rect 51294 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 51914 -3536
rect 51294 -3856 51914 -3772
rect 51294 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 51914 -3856
rect 51294 -7964 51914 -4092
rect 55794 708988 56414 711900
rect 55794 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 56414 708988
rect 55794 708668 56414 708752
rect 55794 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 56414 708668
rect 55794 669454 56414 708432
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4496 56414 20898
rect 55794 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 56414 -4496
rect 55794 -4816 56414 -4732
rect 55794 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 56414 -4816
rect 55794 -7964 56414 -5052
rect 60294 709948 60914 711900
rect 60294 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 60914 709948
rect 60294 709628 60914 709712
rect 60294 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 60914 709628
rect 60294 673954 60914 709392
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5456 60914 25398
rect 60294 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 60914 -5456
rect 60294 -5776 60914 -5692
rect 60294 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 60914 -5776
rect 60294 -7964 60914 -6012
rect 64794 710908 65414 711900
rect 64794 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 65414 710908
rect 64794 710588 65414 710672
rect 64794 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 65414 710588
rect 64794 678454 65414 710352
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6416 65414 29898
rect 64794 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 65414 -6416
rect 64794 -6736 65414 -6652
rect 64794 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 65414 -6736
rect 64794 -7964 65414 -6972
rect 69294 711868 69914 711900
rect 69294 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 69914 711868
rect 69294 711548 69914 711632
rect 69294 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 69914 711548
rect 69294 682954 69914 711312
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7376 69914 34398
rect 69294 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 69914 -7376
rect 69294 -7696 69914 -7612
rect 69294 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 69914 -7696
rect 69294 -7964 69914 -7932
rect 73794 705148 74414 711900
rect 73794 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 74414 705148
rect 73794 704828 74414 704912
rect 73794 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 74414 704828
rect 73794 687454 74414 704592
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 78294 706108 78914 711900
rect 78294 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 78914 706108
rect 78294 705788 78914 705872
rect 78294 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 78914 705788
rect 78294 691954 78914 705552
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 152000 78914 187398
rect 82794 707068 83414 711900
rect 82794 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 83414 707068
rect 82794 706748 83414 706832
rect 82794 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 83414 706748
rect 82794 696454 83414 706512
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 152000 83414 155898
rect 87294 708028 87914 711900
rect 87294 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 87914 708028
rect 87294 707708 87914 707792
rect 87294 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 87914 707708
rect 87294 700954 87914 707472
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 83779 152012 83845 152013
rect 83779 151948 83780 152012
rect 83844 151948 83845 152012
rect 87294 152000 87914 160398
rect 91794 708988 92414 711900
rect 91794 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 92414 708988
rect 91794 708668 92414 708752
rect 91794 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 92414 708668
rect 91794 669454 92414 708432
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 152000 92414 164898
rect 96294 709948 96914 711900
rect 96294 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 96914 709948
rect 96294 709628 96914 709712
rect 96294 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 96914 709628
rect 96294 673954 96914 709392
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 152000 96914 169398
rect 100794 710908 101414 711900
rect 100794 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 101414 710908
rect 100794 710588 101414 710672
rect 100794 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 101414 710588
rect 100794 678454 101414 710352
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 152000 101414 173898
rect 105294 711868 105914 711900
rect 105294 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 105914 711868
rect 105294 711548 105914 711632
rect 105294 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 105914 711548
rect 105294 682954 105914 711312
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 152000 105914 178398
rect 109794 705148 110414 711900
rect 109794 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 110414 705148
rect 109794 704828 110414 704912
rect 109794 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 110414 704828
rect 109794 687454 110414 704592
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 152000 110414 182898
rect 114294 706108 114914 711900
rect 114294 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 114914 706108
rect 114294 705788 114914 705872
rect 114294 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 114914 705788
rect 114294 691954 114914 705552
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 152000 114914 187398
rect 118794 707068 119414 711900
rect 118794 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 119414 707068
rect 118794 706748 119414 706832
rect 118794 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 119414 706748
rect 118794 696454 119414 706512
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 152000 119414 155898
rect 123294 708028 123914 711900
rect 123294 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 123914 708028
rect 123294 707708 123914 707792
rect 123294 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 123914 707708
rect 123294 700954 123914 707472
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122603 152692 122669 152693
rect 122603 152628 122604 152692
rect 122668 152628 122669 152692
rect 122603 152627 122669 152628
rect 83779 151947 83845 151948
rect 82491 151876 82557 151877
rect 82491 151812 82492 151876
rect 82556 151812 82557 151876
rect 82491 151811 82557 151812
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -656 74414 2898
rect 73794 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 74414 -656
rect 73794 -976 74414 -892
rect 73794 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 74414 -976
rect 73794 -7964 74414 -1212
rect 78294 79954 78914 98000
rect 82494 96389 82554 151811
rect 83782 100061 83842 151947
rect 83963 149428 84029 149429
rect 83963 149364 83964 149428
rect 84028 149364 84029 149428
rect 83963 149363 84029 149364
rect 83779 100060 83845 100061
rect 83779 99996 83780 100060
rect 83844 99996 83845 100060
rect 83779 99995 83845 99996
rect 82491 96388 82557 96389
rect 82491 96324 82492 96388
rect 82556 96324 82557 96388
rect 82491 96323 82557 96324
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1616 78914 7398
rect 78294 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 78914 -1616
rect 78294 -1936 78914 -1852
rect 78294 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 78914 -1936
rect 78294 -7964 78914 -2172
rect 82794 84454 83414 98000
rect 83966 97613 84026 149363
rect 84208 147239 84528 147376
rect 84208 147003 84250 147239
rect 84486 147003 84528 147239
rect 84208 146866 84528 147003
rect 114928 147239 115248 147376
rect 114928 147003 114970 147239
rect 115206 147003 115248 147239
rect 114928 146866 115248 147003
rect 99568 115954 99888 115986
rect 99568 115718 99610 115954
rect 99846 115718 99888 115954
rect 99568 115634 99888 115718
rect 99568 115398 99610 115634
rect 99846 115398 99888 115634
rect 99568 115366 99888 115398
rect 84208 111454 84528 111486
rect 84208 111218 84250 111454
rect 84486 111218 84528 111454
rect 84208 111134 84528 111218
rect 84208 110898 84250 111134
rect 84486 110898 84528 111134
rect 84208 110866 84528 110898
rect 114928 111454 115248 111486
rect 114928 111218 114970 111454
rect 115206 111218 115248 111454
rect 114928 111134 115248 111218
rect 114928 110898 114970 111134
rect 115206 110898 115248 111134
rect 114928 110866 115248 110898
rect 122606 109050 122666 152627
rect 123294 152000 123914 160398
rect 127794 708988 128414 711900
rect 127794 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 128414 708988
rect 127794 708668 128414 708752
rect 127794 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 128414 708668
rect 127794 669454 128414 708432
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 124259 152284 124325 152285
rect 124259 152220 124260 152284
rect 124324 152220 124325 152284
rect 124259 152219 124325 152220
rect 122606 108990 123034 109050
rect 99787 100196 99853 100197
rect 99787 100132 99788 100196
rect 99852 100132 99853 100196
rect 99787 100131 99853 100132
rect 84147 99924 84213 99925
rect 84147 99860 84148 99924
rect 84212 99860 84213 99924
rect 84147 99859 84213 99860
rect 85067 99924 85133 99925
rect 85067 99860 85068 99924
rect 85132 99860 85133 99924
rect 85067 99859 85133 99860
rect 86355 99924 86421 99925
rect 86355 99860 86356 99924
rect 86420 99860 86421 99924
rect 86355 99859 86421 99860
rect 89115 99924 89181 99925
rect 89115 99860 89116 99924
rect 89180 99860 89181 99924
rect 89115 99859 89181 99860
rect 90035 99924 90101 99925
rect 90035 99860 90036 99924
rect 90100 99860 90101 99924
rect 90035 99859 90101 99860
rect 90955 99924 91021 99925
rect 90955 99860 90956 99924
rect 91020 99860 91021 99924
rect 93347 99924 93413 99925
rect 93347 99922 93348 99924
rect 90955 99859 91021 99860
rect 93166 99862 93348 99922
rect 83963 97612 84029 97613
rect 83963 97548 83964 97612
rect 84028 97548 84029 97612
rect 83963 97547 84029 97548
rect 84150 89730 84210 99859
rect 85070 99381 85130 99859
rect 85619 99788 85685 99789
rect 85619 99724 85620 99788
rect 85684 99724 85685 99788
rect 85619 99723 85685 99724
rect 85067 99380 85133 99381
rect 85067 99316 85068 99380
rect 85132 99316 85133 99380
rect 85067 99315 85133 99316
rect 84331 98292 84397 98293
rect 84331 98228 84332 98292
rect 84396 98228 84397 98292
rect 84331 98227 84397 98228
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2576 83414 11898
rect 83966 89670 84210 89730
rect 83966 4861 84026 89670
rect 84334 7581 84394 98227
rect 84331 7580 84397 7581
rect 84331 7516 84332 7580
rect 84396 7516 84397 7580
rect 84331 7515 84397 7516
rect 85622 4997 85682 99723
rect 86358 98293 86418 99859
rect 85803 98292 85869 98293
rect 85803 98228 85804 98292
rect 85868 98228 85869 98292
rect 85803 98227 85869 98228
rect 86355 98292 86421 98293
rect 86355 98228 86356 98292
rect 86420 98228 86421 98292
rect 86355 98227 86421 98228
rect 85806 87549 85866 98227
rect 87294 88954 87914 98000
rect 89118 97885 89178 99859
rect 89483 99652 89549 99653
rect 89483 99588 89484 99652
rect 89548 99588 89549 99652
rect 89483 99587 89549 99588
rect 89299 98428 89365 98429
rect 89299 98364 89300 98428
rect 89364 98364 89365 98428
rect 89299 98363 89365 98364
rect 89115 97884 89181 97885
rect 89115 97820 89116 97884
rect 89180 97820 89181 97884
rect 89115 97819 89181 97820
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 85803 87548 85869 87549
rect 85803 87484 85804 87548
rect 85868 87484 85869 87548
rect 85803 87483 85869 87484
rect 87294 52954 87914 88398
rect 89302 88229 89362 98363
rect 89299 88228 89365 88229
rect 89299 88164 89300 88228
rect 89364 88164 89365 88228
rect 89299 88163 89365 88164
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 85619 4996 85685 4997
rect 85619 4932 85620 4996
rect 85684 4932 85685 4996
rect 85619 4931 85685 4932
rect 83963 4860 84029 4861
rect 83963 4796 83964 4860
rect 84028 4796 84029 4860
rect 83963 4795 84029 4796
rect 82794 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 83414 -2576
rect 82794 -2896 83414 -2812
rect 82794 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 83414 -2896
rect 82794 -7964 83414 -3132
rect 87294 -3536 87914 16398
rect 89486 3501 89546 99587
rect 90038 98293 90098 99859
rect 90771 99788 90837 99789
rect 90771 99724 90772 99788
rect 90836 99724 90837 99788
rect 90771 99723 90837 99724
rect 90587 99652 90653 99653
rect 90587 99588 90588 99652
rect 90652 99588 90653 99652
rect 90587 99587 90653 99588
rect 90035 98292 90101 98293
rect 90035 98228 90036 98292
rect 90100 98228 90101 98292
rect 90035 98227 90101 98228
rect 90590 87549 90650 99587
rect 90587 87548 90653 87549
rect 90587 87484 90588 87548
rect 90652 87484 90653 87548
rect 90587 87483 90653 87484
rect 90774 4861 90834 99723
rect 90771 4860 90837 4861
rect 90771 4796 90772 4860
rect 90836 4796 90837 4860
rect 90771 4795 90837 4796
rect 89483 3500 89549 3501
rect 89483 3436 89484 3500
rect 89548 3436 89549 3500
rect 89483 3435 89549 3436
rect 90958 3365 91018 99859
rect 91507 99652 91573 99653
rect 91507 99588 91508 99652
rect 91572 99588 91573 99652
rect 91507 99587 91573 99588
rect 91323 98156 91389 98157
rect 91323 98092 91324 98156
rect 91388 98092 91389 98156
rect 91323 98091 91389 98092
rect 91326 40901 91386 98091
rect 91323 40900 91389 40901
rect 91323 40836 91324 40900
rect 91388 40836 91389 40900
rect 91323 40835 91389 40836
rect 91510 19005 91570 99587
rect 91794 93454 92414 98000
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91507 19004 91573 19005
rect 91507 18940 91508 19004
rect 91572 18940 91573 19004
rect 91507 18939 91573 18940
rect 90955 3364 91021 3365
rect 90955 3300 90956 3364
rect 91020 3300 91021 3364
rect 90955 3299 91021 3300
rect 87294 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 87914 -3536
rect 87294 -3856 87914 -3772
rect 87294 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 87914 -3856
rect 87294 -7964 87914 -4092
rect 91794 -4496 92414 20898
rect 93166 11797 93226 99862
rect 93347 99860 93348 99862
rect 93412 99860 93413 99924
rect 93347 99859 93413 99860
rect 94451 99924 94517 99925
rect 94451 99860 94452 99924
rect 94516 99860 94517 99924
rect 94451 99859 94517 99860
rect 95187 99924 95253 99925
rect 95187 99860 95188 99924
rect 95252 99860 95253 99924
rect 95187 99859 95253 99860
rect 95923 99924 95989 99925
rect 95923 99860 95924 99924
rect 95988 99860 95989 99924
rect 95923 99859 95989 99860
rect 98131 99924 98197 99925
rect 98131 99860 98132 99924
rect 98196 99860 98197 99924
rect 98131 99859 98197 99860
rect 93715 99788 93781 99789
rect 93715 99724 93716 99788
rect 93780 99724 93781 99788
rect 93715 99723 93781 99724
rect 93531 99652 93597 99653
rect 93531 99588 93532 99652
rect 93596 99588 93597 99652
rect 93531 99587 93597 99588
rect 93347 98292 93413 98293
rect 93347 98228 93348 98292
rect 93412 98228 93413 98292
rect 93347 98227 93413 98228
rect 93350 42125 93410 98227
rect 93347 42124 93413 42125
rect 93347 42060 93348 42124
rect 93412 42060 93413 42124
rect 93347 42059 93413 42060
rect 93534 28525 93594 99587
rect 93718 94757 93778 99723
rect 93715 94756 93781 94757
rect 93715 94692 93716 94756
rect 93780 94692 93781 94756
rect 93715 94691 93781 94692
rect 94454 89045 94514 99859
rect 94635 99788 94701 99789
rect 94635 99724 94636 99788
rect 94700 99724 94701 99788
rect 94635 99723 94701 99724
rect 95003 99788 95069 99789
rect 95003 99724 95004 99788
rect 95068 99724 95069 99788
rect 95003 99723 95069 99724
rect 94451 89044 94517 89045
rect 94451 88980 94452 89044
rect 94516 88980 94517 89044
rect 94451 88979 94517 88980
rect 94638 40765 94698 99723
rect 94819 97884 94885 97885
rect 94819 97820 94820 97884
rect 94884 97820 94885 97884
rect 94819 97819 94885 97820
rect 94635 40764 94701 40765
rect 94635 40700 94636 40764
rect 94700 40700 94701 40764
rect 94635 40699 94701 40700
rect 94822 36413 94882 97819
rect 94819 36412 94885 36413
rect 94819 36348 94820 36412
rect 94884 36348 94885 36412
rect 94819 36347 94885 36348
rect 93531 28524 93597 28525
rect 93531 28460 93532 28524
rect 93596 28460 93597 28524
rect 93531 28459 93597 28460
rect 95006 20093 95066 99723
rect 95190 98293 95250 99859
rect 95187 98292 95253 98293
rect 95187 98228 95188 98292
rect 95252 98228 95253 98292
rect 95187 98227 95253 98228
rect 95739 97612 95805 97613
rect 95739 97548 95740 97612
rect 95804 97548 95805 97612
rect 95739 97547 95805 97548
rect 95742 40629 95802 97547
rect 95739 40628 95805 40629
rect 95739 40564 95740 40628
rect 95804 40564 95805 40628
rect 95739 40563 95805 40564
rect 95926 37229 95986 99859
rect 96107 99788 96173 99789
rect 96107 99724 96108 99788
rect 96172 99724 96173 99788
rect 96107 99723 96173 99724
rect 97763 99788 97829 99789
rect 97763 99724 97764 99788
rect 97828 99724 97829 99788
rect 97763 99723 97829 99724
rect 95923 37228 95989 37229
rect 95923 37164 95924 37228
rect 95988 37164 95989 37228
rect 95923 37163 95989 37164
rect 95003 20092 95069 20093
rect 95003 20028 95004 20092
rect 95068 20028 95069 20092
rect 95003 20027 95069 20028
rect 93163 11796 93229 11797
rect 93163 11732 93164 11796
rect 93228 11732 93229 11796
rect 93163 11731 93229 11732
rect 96110 7581 96170 99723
rect 96294 97954 96914 98000
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 97579 97612 97645 97613
rect 97579 97548 97580 97612
rect 97644 97548 97645 97612
rect 97579 97547 97645 97548
rect 97395 97476 97461 97477
rect 97395 97412 97396 97476
rect 97460 97412 97461 97476
rect 97395 97411 97461 97412
rect 96294 61954 96914 97398
rect 97211 97204 97277 97205
rect 97211 97140 97212 97204
rect 97276 97140 97277 97204
rect 97211 97139 97277 97140
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 97214 38317 97274 97139
rect 97211 38316 97277 38317
rect 97211 38252 97212 38316
rect 97276 38252 97277 38316
rect 97211 38251 97277 38252
rect 97398 37093 97458 97411
rect 97395 37092 97461 37093
rect 97395 37028 97396 37092
rect 97460 37028 97461 37092
rect 97395 37027 97461 37028
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96107 7580 96173 7581
rect 96107 7516 96108 7580
rect 96172 7516 96173 7580
rect 96107 7515 96173 7516
rect 91794 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 92414 -4496
rect 91794 -4816 92414 -4732
rect 91794 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 92414 -4816
rect 91794 -7964 92414 -5052
rect 96294 -5456 96914 25398
rect 97582 9349 97642 97547
rect 97766 9485 97826 99723
rect 98134 97613 98194 99859
rect 99790 99789 99850 100131
rect 110643 100060 110709 100061
rect 110643 99996 110644 100060
rect 110708 99996 110709 100060
rect 110643 99995 110709 99996
rect 100523 99924 100589 99925
rect 100523 99860 100524 99924
rect 100588 99860 100589 99924
rect 100523 99859 100589 99860
rect 101811 99924 101877 99925
rect 101811 99860 101812 99924
rect 101876 99860 101877 99924
rect 101811 99859 101877 99860
rect 102179 99924 102245 99925
rect 102179 99860 102180 99924
rect 102244 99860 102245 99924
rect 102179 99859 102245 99860
rect 102915 99924 102981 99925
rect 102915 99860 102916 99924
rect 102980 99860 102981 99924
rect 102915 99859 102981 99860
rect 105307 99924 105373 99925
rect 105307 99860 105308 99924
rect 105372 99860 105373 99924
rect 105307 99859 105373 99860
rect 106043 99924 106109 99925
rect 106043 99860 106044 99924
rect 106108 99860 106109 99924
rect 106043 99859 106109 99860
rect 107331 99924 107397 99925
rect 107331 99860 107332 99924
rect 107396 99860 107397 99924
rect 107331 99859 107397 99860
rect 108251 99924 108317 99925
rect 108251 99860 108252 99924
rect 108316 99860 108317 99924
rect 108251 99859 108317 99860
rect 109907 99924 109973 99925
rect 109907 99860 109908 99924
rect 109972 99922 109973 99924
rect 109972 99862 110154 99922
rect 109972 99860 109973 99862
rect 109907 99859 109973 99860
rect 99787 99788 99853 99789
rect 99787 99724 99788 99788
rect 99852 99724 99853 99788
rect 99787 99723 99853 99724
rect 98683 99516 98749 99517
rect 98683 99452 98684 99516
rect 98748 99452 98749 99516
rect 98683 99451 98749 99452
rect 98131 97612 98197 97613
rect 98131 97548 98132 97612
rect 98196 97548 98197 97612
rect 98131 97547 98197 97548
rect 98686 38181 98746 99451
rect 98867 97612 98933 97613
rect 98867 97548 98868 97612
rect 98932 97548 98933 97612
rect 98867 97547 98933 97548
rect 99235 97612 99301 97613
rect 99235 97548 99236 97612
rect 99300 97548 99301 97612
rect 99235 97547 99301 97548
rect 98683 38180 98749 38181
rect 98683 38116 98684 38180
rect 98748 38116 98749 38180
rect 98683 38115 98749 38116
rect 98870 24445 98930 97547
rect 99051 97476 99117 97477
rect 99051 97412 99052 97476
rect 99116 97412 99117 97476
rect 99051 97411 99117 97412
rect 98867 24444 98933 24445
rect 98867 24380 98868 24444
rect 98932 24380 98933 24444
rect 98867 24379 98933 24380
rect 99054 21453 99114 97411
rect 99051 21452 99117 21453
rect 99051 21388 99052 21452
rect 99116 21388 99117 21452
rect 99051 21387 99117 21388
rect 97763 9484 97829 9485
rect 97763 9420 97764 9484
rect 97828 9420 97829 9484
rect 97763 9419 97829 9420
rect 97579 9348 97645 9349
rect 97579 9284 97580 9348
rect 97644 9284 97645 9348
rect 97579 9283 97645 9284
rect 99238 6629 99298 97547
rect 99790 97069 99850 99723
rect 100155 98428 100221 98429
rect 100155 98364 100156 98428
rect 100220 98364 100221 98428
rect 100155 98363 100221 98364
rect 99971 98292 100037 98293
rect 99971 98228 99972 98292
rect 100036 98228 100037 98292
rect 99971 98227 100037 98228
rect 99787 97068 99853 97069
rect 99787 97004 99788 97068
rect 99852 97004 99853 97068
rect 99787 97003 99853 97004
rect 99974 9213 100034 98227
rect 100158 27165 100218 98363
rect 100339 98156 100405 98157
rect 100339 98092 100340 98156
rect 100404 98092 100405 98156
rect 100339 98091 100405 98092
rect 100155 27164 100221 27165
rect 100155 27100 100156 27164
rect 100220 27100 100221 27164
rect 100155 27099 100221 27100
rect 99971 9212 100037 9213
rect 99971 9148 99972 9212
rect 100036 9148 100037 9212
rect 99971 9147 100037 9148
rect 100342 9077 100402 98091
rect 100526 94621 100586 99859
rect 101627 99516 101693 99517
rect 101627 99452 101628 99516
rect 101692 99452 101693 99516
rect 101627 99451 101693 99452
rect 100523 94620 100589 94621
rect 100523 94556 100524 94620
rect 100588 94556 100589 94620
rect 100523 94555 100589 94556
rect 100794 66454 101414 98000
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100339 9076 100405 9077
rect 100339 9012 100340 9076
rect 100404 9012 100405 9076
rect 100339 9011 100405 9012
rect 99235 6628 99301 6629
rect 99235 6564 99236 6628
rect 99300 6564 99301 6628
rect 99235 6563 99301 6564
rect 96294 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 96914 -5456
rect 96294 -5776 96914 -5692
rect 96294 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 96914 -5776
rect 96294 -7964 96914 -6012
rect 100794 -6416 101414 29898
rect 101630 25533 101690 99451
rect 101814 98293 101874 99859
rect 102182 98293 102242 99859
rect 102918 98293 102978 99859
rect 103283 99788 103349 99789
rect 103283 99724 103284 99788
rect 103348 99724 103349 99788
rect 103283 99723 103349 99724
rect 103099 99652 103165 99653
rect 103099 99588 103100 99652
rect 103164 99588 103165 99652
rect 103099 99587 103165 99588
rect 101811 98292 101877 98293
rect 101811 98228 101812 98292
rect 101876 98228 101877 98292
rect 101811 98227 101877 98228
rect 102179 98292 102245 98293
rect 102179 98228 102180 98292
rect 102244 98228 102245 98292
rect 102179 98227 102245 98228
rect 102915 98292 102981 98293
rect 102915 98228 102916 98292
rect 102980 98228 102981 98292
rect 102915 98227 102981 98228
rect 101995 95708 102061 95709
rect 101995 95644 101996 95708
rect 102060 95644 102061 95708
rect 101995 95643 102061 95644
rect 101811 95572 101877 95573
rect 101811 95508 101812 95572
rect 101876 95508 101877 95572
rect 101811 95507 101877 95508
rect 101627 25532 101693 25533
rect 101627 25468 101628 25532
rect 101692 25468 101693 25532
rect 101627 25467 101693 25468
rect 101814 22949 101874 95507
rect 101811 22948 101877 22949
rect 101811 22884 101812 22948
rect 101876 22884 101877 22948
rect 101811 22883 101877 22884
rect 101998 8941 102058 95643
rect 102915 95572 102981 95573
rect 102915 95508 102916 95572
rect 102980 95508 102981 95572
rect 102915 95507 102981 95508
rect 102731 91764 102797 91765
rect 102731 91700 102732 91764
rect 102796 91700 102797 91764
rect 102731 91699 102797 91700
rect 102734 84965 102794 91699
rect 102731 84964 102797 84965
rect 102731 84900 102732 84964
rect 102796 84900 102797 84964
rect 102731 84899 102797 84900
rect 102918 27029 102978 95507
rect 102915 27028 102981 27029
rect 102915 26964 102916 27028
rect 102980 26964 102981 27028
rect 102915 26963 102981 26964
rect 103102 26893 103162 99587
rect 103099 26892 103165 26893
rect 103099 26828 103100 26892
rect 103164 26828 103165 26892
rect 103099 26827 103165 26828
rect 103286 10437 103346 99723
rect 105310 98293 105370 99859
rect 103651 98292 103717 98293
rect 103651 98228 103652 98292
rect 103716 98228 103717 98292
rect 103651 98227 103717 98228
rect 105307 98292 105373 98293
rect 105307 98228 105308 98292
rect 105372 98228 105373 98292
rect 105307 98227 105373 98228
rect 103654 95573 103714 98227
rect 104203 96524 104269 96525
rect 104203 96460 104204 96524
rect 104268 96460 104269 96524
rect 104203 96459 104269 96460
rect 103651 95572 103717 95573
rect 103651 95508 103652 95572
rect 103716 95508 103717 95572
rect 103651 95507 103717 95508
rect 103283 10436 103349 10437
rect 103283 10372 103284 10436
rect 103348 10372 103349 10436
rect 103283 10371 103349 10372
rect 104206 10301 104266 96459
rect 105123 96252 105189 96253
rect 105123 96188 105124 96252
rect 105188 96188 105189 96252
rect 105123 96187 105189 96188
rect 104571 95708 104637 95709
rect 104571 95644 104572 95708
rect 104636 95644 104637 95708
rect 104571 95643 104637 95644
rect 104387 95572 104453 95573
rect 104387 95508 104388 95572
rect 104452 95508 104453 95572
rect 104387 95507 104453 95508
rect 104390 28253 104450 95507
rect 104574 28389 104634 95643
rect 105126 29613 105186 96187
rect 105294 70954 105914 98000
rect 106046 84829 106106 99859
rect 107147 96388 107213 96389
rect 107147 96324 107148 96388
rect 107212 96324 107213 96388
rect 107147 96323 107213 96324
rect 106963 96252 107029 96253
rect 106963 96188 106964 96252
rect 107028 96188 107029 96252
rect 106963 96187 107029 96188
rect 106043 84828 106109 84829
rect 106043 84764 106044 84828
rect 106108 84764 106109 84828
rect 106043 84763 106109 84764
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105123 29612 105189 29613
rect 105123 29548 105124 29612
rect 105188 29548 105189 29612
rect 105123 29547 105189 29548
rect 104571 28388 104637 28389
rect 104571 28324 104572 28388
rect 104636 28324 104637 28388
rect 104571 28323 104637 28324
rect 104387 28252 104453 28253
rect 104387 28188 104388 28252
rect 104452 28188 104453 28252
rect 104387 28187 104453 28188
rect 104203 10300 104269 10301
rect 104203 10236 104204 10300
rect 104268 10236 104269 10300
rect 104203 10235 104269 10236
rect 101995 8940 102061 8941
rect 101995 8876 101996 8940
rect 102060 8876 102061 8940
rect 101995 8875 102061 8876
rect 100794 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 101414 -6416
rect 100794 -6736 101414 -6652
rect 100794 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 101414 -6736
rect 100794 -7964 101414 -6972
rect 105294 -7376 105914 34398
rect 106966 30973 107026 96187
rect 107150 31109 107210 96323
rect 107147 31108 107213 31109
rect 107147 31044 107148 31108
rect 107212 31044 107213 31108
rect 107147 31043 107213 31044
rect 106963 30972 107029 30973
rect 106963 30908 106964 30972
rect 107028 30908 107029 30972
rect 106963 30907 107029 30908
rect 107334 13293 107394 99859
rect 108067 99788 108133 99789
rect 108067 99724 108068 99788
rect 108132 99724 108133 99788
rect 108067 99723 108133 99724
rect 107515 99652 107581 99653
rect 107515 99588 107516 99652
rect 107580 99588 107581 99652
rect 107515 99587 107581 99588
rect 107331 13292 107397 13293
rect 107331 13228 107332 13292
rect 107396 13228 107397 13292
rect 107331 13227 107397 13228
rect 107518 11661 107578 99587
rect 108070 95437 108130 99723
rect 108254 99653 108314 99859
rect 108251 99652 108317 99653
rect 108251 99588 108252 99652
rect 108316 99588 108317 99652
rect 108251 99587 108317 99588
rect 108435 99652 108501 99653
rect 108435 99588 108436 99652
rect 108500 99588 108501 99652
rect 108435 99587 108501 99588
rect 108067 95436 108133 95437
rect 108067 95372 108068 95436
rect 108132 95372 108133 95436
rect 108067 95371 108133 95372
rect 108438 39405 108498 99587
rect 110094 98157 110154 99862
rect 110091 98156 110157 98157
rect 110091 98092 110092 98156
rect 110156 98092 110157 98156
rect 110091 98091 110157 98092
rect 109355 96796 109421 96797
rect 109355 96732 109356 96796
rect 109420 96732 109421 96796
rect 109355 96731 109421 96732
rect 108803 96660 108869 96661
rect 108803 96596 108804 96660
rect 108868 96596 108869 96660
rect 108803 96595 108869 96596
rect 108619 96252 108685 96253
rect 108619 96188 108620 96252
rect 108684 96188 108685 96252
rect 108619 96187 108685 96188
rect 108435 39404 108501 39405
rect 108435 39340 108436 39404
rect 108500 39340 108501 39404
rect 108435 39339 108501 39340
rect 108622 24309 108682 96187
rect 108619 24308 108685 24309
rect 108619 24244 108620 24308
rect 108684 24244 108685 24308
rect 108619 24243 108685 24244
rect 108806 13157 108866 96595
rect 109358 24173 109418 96731
rect 109539 96252 109605 96253
rect 109539 96188 109540 96252
rect 109604 96188 109605 96252
rect 109539 96187 109605 96188
rect 109355 24172 109421 24173
rect 109355 24108 109356 24172
rect 109420 24108 109421 24172
rect 109355 24107 109421 24108
rect 108803 13156 108869 13157
rect 108803 13092 108804 13156
rect 108868 13092 108869 13156
rect 108803 13091 108869 13092
rect 109542 13021 109602 96187
rect 109794 75454 110414 98000
rect 110646 93533 110706 99995
rect 111011 99924 111077 99925
rect 111011 99860 111012 99924
rect 111076 99860 111077 99924
rect 111011 99859 111077 99860
rect 111563 99924 111629 99925
rect 111563 99860 111564 99924
rect 111628 99860 111629 99924
rect 111563 99859 111629 99860
rect 116347 99924 116413 99925
rect 116347 99860 116348 99924
rect 116412 99860 116413 99924
rect 116347 99859 116413 99860
rect 117083 99924 117149 99925
rect 117083 99860 117084 99924
rect 117148 99860 117149 99924
rect 117083 99859 117149 99860
rect 117819 99924 117885 99925
rect 117819 99860 117820 99924
rect 117884 99860 117885 99924
rect 117819 99859 117885 99860
rect 120763 99924 120829 99925
rect 120763 99860 120764 99924
rect 120828 99860 120829 99924
rect 120763 99859 120829 99860
rect 111014 96525 111074 99859
rect 111195 99380 111261 99381
rect 111195 99316 111196 99380
rect 111260 99316 111261 99380
rect 111195 99315 111261 99316
rect 111011 96524 111077 96525
rect 111011 96460 111012 96524
rect 111076 96460 111077 96524
rect 111011 96459 111077 96460
rect 111011 96388 111077 96389
rect 111011 96324 111012 96388
rect 111076 96324 111077 96388
rect 111011 96323 111077 96324
rect 110643 93532 110709 93533
rect 110643 93468 110644 93532
rect 110708 93468 110709 93532
rect 110643 93467 110709 93468
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109539 13020 109605 13021
rect 109539 12956 109540 13020
rect 109604 12956 109605 13020
rect 109539 12955 109605 12956
rect 107515 11660 107581 11661
rect 107515 11596 107516 11660
rect 107580 11596 107581 11660
rect 107515 11595 107581 11596
rect 105294 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 105914 -7376
rect 105294 -7696 105914 -7612
rect 105294 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 105914 -7696
rect 105294 -7964 105914 -7932
rect 109794 3454 110414 38898
rect 111014 14789 111074 96323
rect 111198 36957 111258 99315
rect 111379 95572 111445 95573
rect 111379 95508 111380 95572
rect 111444 95508 111445 95572
rect 111379 95507 111445 95508
rect 111195 36956 111261 36957
rect 111195 36892 111196 36956
rect 111260 36892 111261 36956
rect 111195 36891 111261 36892
rect 111382 14925 111442 95507
rect 111566 93261 111626 99859
rect 114139 99788 114205 99789
rect 114139 99724 114140 99788
rect 114204 99724 114205 99788
rect 114139 99723 114205 99724
rect 112483 97068 112549 97069
rect 112483 97004 112484 97068
rect 112548 97004 112549 97068
rect 112483 97003 112549 97004
rect 111563 93260 111629 93261
rect 111563 93196 111564 93260
rect 111628 93196 111629 93260
rect 111563 93195 111629 93196
rect 112486 93125 112546 97003
rect 113035 96932 113101 96933
rect 113035 96868 113036 96932
rect 113100 96868 113101 96932
rect 113035 96867 113101 96868
rect 113587 96932 113653 96933
rect 113587 96868 113588 96932
rect 113652 96868 113653 96932
rect 113587 96867 113653 96868
rect 112667 96796 112733 96797
rect 112667 96732 112668 96796
rect 112732 96732 112733 96796
rect 112667 96731 112733 96732
rect 112483 93124 112549 93125
rect 112483 93060 112484 93124
rect 112548 93060 112549 93124
rect 112483 93059 112549 93060
rect 112670 36821 112730 96731
rect 112851 96660 112917 96661
rect 112851 96596 112852 96660
rect 112916 96596 112917 96660
rect 112851 96595 112917 96596
rect 112667 36820 112733 36821
rect 112667 36756 112668 36820
rect 112732 36756 112733 36820
rect 112667 36755 112733 36756
rect 111379 14924 111445 14925
rect 111379 14860 111380 14924
rect 111444 14860 111445 14924
rect 111379 14859 111445 14860
rect 111011 14788 111077 14789
rect 111011 14724 111012 14788
rect 111076 14724 111077 14788
rect 111011 14723 111077 14724
rect 112854 14517 112914 96595
rect 113038 14653 113098 96867
rect 113590 33829 113650 96867
rect 113955 96796 114021 96797
rect 113955 96732 113956 96796
rect 114020 96732 114021 96796
rect 113955 96731 114021 96732
rect 113771 96660 113837 96661
rect 113771 96596 113772 96660
rect 113836 96596 113837 96660
rect 113771 96595 113837 96596
rect 113587 33828 113653 33829
rect 113587 33764 113588 33828
rect 113652 33764 113653 33828
rect 113587 33763 113653 33764
rect 113774 32605 113834 96595
rect 113771 32604 113837 32605
rect 113771 32540 113772 32604
rect 113836 32540 113837 32604
rect 113771 32539 113837 32540
rect 113958 16149 114018 96731
rect 113955 16148 114021 16149
rect 113955 16084 113956 16148
rect 114020 16084 114021 16148
rect 113955 16083 114021 16084
rect 114142 16013 114202 99723
rect 114294 79954 114914 98000
rect 116350 96933 116410 99859
rect 116715 99652 116781 99653
rect 116715 99588 116716 99652
rect 116780 99588 116781 99652
rect 116715 99587 116781 99588
rect 116347 96932 116413 96933
rect 116347 96868 116348 96932
rect 116412 96868 116413 96932
rect 116347 96867 116413 96868
rect 115611 96796 115677 96797
rect 115611 96732 115612 96796
rect 115676 96732 115677 96796
rect 115611 96731 115677 96732
rect 115614 90813 115674 96731
rect 115795 96660 115861 96661
rect 115795 96596 115796 96660
rect 115860 96596 115861 96660
rect 115795 96595 115861 96596
rect 115611 90812 115677 90813
rect 115611 90748 115612 90812
rect 115676 90748 115677 90812
rect 115611 90747 115677 90748
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114139 16012 114205 16013
rect 114139 15948 114140 16012
rect 114204 15948 114205 16012
rect 114139 15947 114205 15948
rect 113035 14652 113101 14653
rect 113035 14588 113036 14652
rect 113100 14588 113101 14652
rect 113035 14587 113101 14588
rect 112851 14516 112917 14517
rect 112851 14452 112852 14516
rect 112916 14452 112917 14516
rect 112851 14451 112917 14452
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -656 110414 2898
rect 109794 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 110414 -656
rect 109794 -976 110414 -892
rect 109794 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 110414 -976
rect 109794 -7964 110414 -1212
rect 114294 7954 114914 43398
rect 115798 15877 115858 96595
rect 116718 38045 116778 99587
rect 116899 97476 116965 97477
rect 116899 97412 116900 97476
rect 116964 97412 116965 97476
rect 116899 97411 116965 97412
rect 116715 38044 116781 38045
rect 116715 37980 116716 38044
rect 116780 37980 116781 38044
rect 116715 37979 116781 37980
rect 116902 35733 116962 97411
rect 116899 35732 116965 35733
rect 116899 35668 116900 35732
rect 116964 35668 116965 35732
rect 116899 35667 116965 35668
rect 117086 35597 117146 99859
rect 117267 99516 117333 99517
rect 117267 99452 117268 99516
rect 117332 99452 117333 99516
rect 117267 99451 117333 99452
rect 117270 90677 117330 99451
rect 117267 90676 117333 90677
rect 117267 90612 117268 90676
rect 117332 90612 117333 90676
rect 117267 90611 117333 90612
rect 117822 37909 117882 99859
rect 118187 99788 118253 99789
rect 118187 99724 118188 99788
rect 118252 99724 118253 99788
rect 118187 99723 118253 99724
rect 119659 99788 119725 99789
rect 119659 99724 119660 99788
rect 119724 99724 119725 99788
rect 119659 99723 119725 99724
rect 118003 99652 118069 99653
rect 118003 99588 118004 99652
rect 118068 99588 118069 99652
rect 118003 99587 118069 99588
rect 117819 37908 117885 37909
rect 117819 37844 117820 37908
rect 117884 37844 117885 37908
rect 117819 37843 117885 37844
rect 117083 35596 117149 35597
rect 117083 35532 117084 35596
rect 117148 35532 117149 35596
rect 117083 35531 117149 35532
rect 118006 35325 118066 99587
rect 118190 35461 118250 99723
rect 118555 97204 118621 97205
rect 118555 97140 118556 97204
rect 118620 97140 118621 97204
rect 118555 97139 118621 97140
rect 118371 97068 118437 97069
rect 118371 97004 118372 97068
rect 118436 97004 118437 97068
rect 118371 97003 118437 97004
rect 118187 35460 118253 35461
rect 118187 35396 118188 35460
rect 118252 35396 118253 35460
rect 118187 35395 118253 35396
rect 118003 35324 118069 35325
rect 118003 35260 118004 35324
rect 118068 35260 118069 35324
rect 118003 35259 118069 35260
rect 118374 17509 118434 97003
rect 118371 17508 118437 17509
rect 118371 17444 118372 17508
rect 118436 17444 118437 17508
rect 118371 17443 118437 17444
rect 118558 17373 118618 97139
rect 118794 84454 119414 98000
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118555 17372 118621 17373
rect 118555 17308 118556 17372
rect 118620 17308 118621 17372
rect 118555 17307 118621 17308
rect 115795 15876 115861 15877
rect 115795 15812 115796 15876
rect 115860 15812 115861 15876
rect 115795 15811 115861 15812
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1616 114914 7398
rect 114294 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 114914 -1616
rect 114294 -1936 114914 -1852
rect 114294 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 114914 -1936
rect 114294 -7964 114914 -2172
rect 118794 12454 119414 47898
rect 119662 32469 119722 99723
rect 119843 97204 119909 97205
rect 119843 97140 119844 97204
rect 119908 97140 119909 97204
rect 119843 97139 119909 97140
rect 120579 97204 120645 97205
rect 120579 97140 120580 97204
rect 120644 97140 120645 97204
rect 120579 97139 120645 97140
rect 119659 32468 119725 32469
rect 119659 32404 119660 32468
rect 119724 32404 119725 32468
rect 119659 32403 119725 32404
rect 119846 18869 119906 97139
rect 120582 90541 120642 97139
rect 120766 97069 120826 99859
rect 120947 99788 121013 99789
rect 120947 99724 120948 99788
rect 121012 99724 121013 99788
rect 120947 99723 121013 99724
rect 122419 99788 122485 99789
rect 122419 99724 122420 99788
rect 122484 99724 122485 99788
rect 122419 99723 122485 99724
rect 122603 99788 122669 99789
rect 122603 99724 122604 99788
rect 122668 99724 122669 99788
rect 122603 99723 122669 99724
rect 120763 97068 120829 97069
rect 120763 97004 120764 97068
rect 120828 97004 120829 97068
rect 120763 97003 120829 97004
rect 120763 96932 120829 96933
rect 120763 96868 120764 96932
rect 120828 96868 120829 96932
rect 120763 96867 120829 96868
rect 120579 90540 120645 90541
rect 120579 90476 120580 90540
rect 120644 90476 120645 90540
rect 120579 90475 120645 90476
rect 119843 18868 119909 18869
rect 119843 18804 119844 18868
rect 119908 18804 119909 18868
rect 119843 18803 119909 18804
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2576 119414 11898
rect 120766 6357 120826 96867
rect 120950 35189 121010 99723
rect 122051 98428 122117 98429
rect 122051 98364 122052 98428
rect 122116 98364 122117 98428
rect 122051 98363 122117 98364
rect 121131 97340 121197 97341
rect 121131 97276 121132 97340
rect 121196 97276 121197 97340
rect 121131 97275 121197 97276
rect 120947 35188 121013 35189
rect 120947 35124 120948 35188
rect 121012 35124 121013 35188
rect 120947 35123 121013 35124
rect 121134 6493 121194 97275
rect 121131 6492 121197 6493
rect 121131 6428 121132 6492
rect 121196 6428 121197 6492
rect 121131 6427 121197 6428
rect 120763 6356 120829 6357
rect 120763 6292 120764 6356
rect 120828 6292 120829 6356
rect 120763 6291 120829 6292
rect 122054 6221 122114 98363
rect 122235 96796 122301 96797
rect 122235 96732 122236 96796
rect 122300 96732 122301 96796
rect 122235 96731 122301 96732
rect 122238 18733 122298 96731
rect 122235 18732 122301 18733
rect 122235 18668 122236 18732
rect 122300 18668 122301 18732
rect 122235 18667 122301 18668
rect 122422 17237 122482 99723
rect 122606 90405 122666 99723
rect 122787 98292 122853 98293
rect 122787 98228 122788 98292
rect 122852 98228 122853 98292
rect 122787 98227 122853 98228
rect 122790 95845 122850 98227
rect 122974 97749 123034 108990
rect 124075 99924 124141 99925
rect 124075 99860 124076 99924
rect 124140 99860 124141 99924
rect 124075 99859 124141 99860
rect 122971 97748 123037 97749
rect 122971 97684 122972 97748
rect 123036 97684 123037 97748
rect 122971 97683 123037 97684
rect 122971 97612 123037 97613
rect 122971 97548 122972 97612
rect 123036 97548 123037 97612
rect 122971 97547 123037 97548
rect 122787 95844 122853 95845
rect 122787 95780 122788 95844
rect 122852 95780 122853 95844
rect 122787 95779 122853 95780
rect 122603 90404 122669 90405
rect 122603 90340 122604 90404
rect 122668 90340 122669 90404
rect 122603 90339 122669 90340
rect 122974 21317 123034 97547
rect 123294 88954 123914 98000
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 122971 21316 123037 21317
rect 122971 21252 122972 21316
rect 123036 21252 123037 21316
rect 122971 21251 123037 21252
rect 122419 17236 122485 17237
rect 122419 17172 122420 17236
rect 122484 17172 122485 17236
rect 122419 17171 122485 17172
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 122051 6220 122117 6221
rect 122051 6156 122052 6220
rect 122116 6156 122117 6220
rect 122051 6155 122117 6156
rect 118794 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 119414 -2576
rect 118794 -2896 119414 -2812
rect 118794 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 119414 -2896
rect 118794 -7964 119414 -3132
rect 123294 -3536 123914 16398
rect 124078 4861 124138 99859
rect 124262 92445 124322 152219
rect 124443 152012 124509 152013
rect 124443 151948 124444 152012
rect 124508 151948 124509 152012
rect 127794 152000 128414 164898
rect 132294 709948 132914 711900
rect 132294 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 132914 709948
rect 132294 709628 132914 709712
rect 132294 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 132914 709628
rect 132294 673954 132914 709392
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 124443 151947 124509 151948
rect 124446 100197 124506 151947
rect 128859 150516 128925 150517
rect 128859 150452 128860 150516
rect 128924 150452 128925 150516
rect 128859 150451 128925 150452
rect 124443 100196 124509 100197
rect 124443 100132 124444 100196
rect 124508 100132 124509 100196
rect 124443 100131 124509 100132
rect 124811 99924 124877 99925
rect 124811 99860 124812 99924
rect 124876 99860 124877 99924
rect 124811 99859 124877 99860
rect 126099 99924 126165 99925
rect 126099 99860 126100 99924
rect 126164 99860 126165 99924
rect 126099 99859 126165 99860
rect 126651 99924 126717 99925
rect 126651 99860 126652 99924
rect 126716 99860 126717 99924
rect 126651 99859 126717 99860
rect 124259 92444 124325 92445
rect 124259 92380 124260 92444
rect 124324 92380 124325 92444
rect 124259 92379 124325 92380
rect 124814 79389 124874 99859
rect 126102 98293 126162 99859
rect 126654 98970 126714 99859
rect 126286 98910 126714 98970
rect 126099 98292 126165 98293
rect 126099 98228 126100 98292
rect 126164 98228 126165 98292
rect 126099 98227 126165 98228
rect 124995 97068 125061 97069
rect 124995 97004 124996 97068
rect 125060 97004 125061 97068
rect 124995 97003 125061 97004
rect 124811 79388 124877 79389
rect 124811 79324 124812 79388
rect 124876 79324 124877 79388
rect 124811 79323 124877 79324
rect 124998 36685 125058 97003
rect 125363 96796 125429 96797
rect 125363 96732 125364 96796
rect 125428 96732 125429 96796
rect 125363 96731 125429 96732
rect 125179 96660 125245 96661
rect 125179 96596 125180 96660
rect 125244 96596 125245 96660
rect 125179 96595 125245 96596
rect 124995 36684 125061 36685
rect 124995 36620 124996 36684
rect 125060 36620 125061 36684
rect 124995 36619 125061 36620
rect 125182 22813 125242 96595
rect 125179 22812 125245 22813
rect 125179 22748 125180 22812
rect 125244 22748 125245 22812
rect 125179 22747 125245 22748
rect 125366 18597 125426 96731
rect 126286 39269 126346 98910
rect 126467 98292 126533 98293
rect 126467 98228 126468 98292
rect 126532 98228 126533 98292
rect 126467 98227 126533 98228
rect 126283 39268 126349 39269
rect 126283 39204 126284 39268
rect 126348 39204 126349 39268
rect 126283 39203 126349 39204
rect 126470 36549 126530 98227
rect 126651 98156 126717 98157
rect 126651 98092 126652 98156
rect 126716 98092 126717 98156
rect 126651 98091 126717 98092
rect 126467 36548 126533 36549
rect 126467 36484 126468 36548
rect 126532 36484 126533 36548
rect 126467 36483 126533 36484
rect 126654 22677 126714 98091
rect 126835 97340 126901 97341
rect 126835 97276 126836 97340
rect 126900 97276 126901 97340
rect 126835 97275 126901 97276
rect 126651 22676 126717 22677
rect 126651 22612 126652 22676
rect 126716 22612 126717 22676
rect 126651 22611 126717 22612
rect 126838 19957 126898 97275
rect 127794 93454 128414 98000
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 128862 38725 128922 150451
rect 132294 133954 132914 169398
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 128859 38724 128925 38725
rect 128859 38660 128860 38724
rect 128924 38660 128925 38724
rect 128859 38659 128925 38660
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 126835 19956 126901 19957
rect 126835 19892 126836 19956
rect 126900 19892 126901 19956
rect 126835 19891 126901 19892
rect 125363 18596 125429 18597
rect 125363 18532 125364 18596
rect 125428 18532 125429 18596
rect 125363 18531 125429 18532
rect 124075 4860 124141 4861
rect 124075 4796 124076 4860
rect 124140 4796 124141 4860
rect 124075 4795 124141 4796
rect 123294 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 123914 -3536
rect 123294 -3856 123914 -3772
rect 123294 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 123914 -3856
rect 123294 -7964 123914 -4092
rect 127794 -4496 128414 20898
rect 127794 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 128414 -4496
rect 127794 -4816 128414 -4732
rect 127794 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 128414 -4816
rect 127794 -7964 128414 -5052
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5456 132914 25398
rect 132294 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 132914 -5456
rect 132294 -5776 132914 -5692
rect 132294 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 132914 -5776
rect 132294 -7964 132914 -6012
rect 136794 710908 137414 711900
rect 136794 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 137414 710908
rect 136794 710588 137414 710672
rect 136794 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 137414 710588
rect 136794 678454 137414 710352
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 138454 137414 173898
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6416 137414 29898
rect 136794 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 137414 -6416
rect 136794 -6736 137414 -6652
rect 136794 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 137414 -6736
rect 136794 -7964 137414 -6972
rect 141294 711868 141914 711900
rect 141294 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 141914 711868
rect 141294 711548 141914 711632
rect 141294 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 141914 711548
rect 141294 682954 141914 711312
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7376 141914 34398
rect 141294 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 141914 -7376
rect 141294 -7696 141914 -7612
rect 141294 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 141914 -7696
rect 141294 -7964 141914 -7932
rect 145794 705148 146414 711900
rect 145794 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 146414 705148
rect 145794 704828 146414 704912
rect 145794 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 146414 704828
rect 145794 687454 146414 704592
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -656 146414 2898
rect 145794 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 146414 -656
rect 145794 -976 146414 -892
rect 145794 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 146414 -976
rect 145794 -7964 146414 -1212
rect 150294 706108 150914 711900
rect 150294 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 150914 706108
rect 150294 705788 150914 705872
rect 150294 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 150914 705788
rect 150294 691954 150914 705552
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1616 150914 7398
rect 150294 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 150914 -1616
rect 150294 -1936 150914 -1852
rect 150294 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 150914 -1936
rect 150294 -7964 150914 -2172
rect 154794 707068 155414 711900
rect 154794 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 155414 707068
rect 154794 706748 155414 706832
rect 154794 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 155414 706748
rect 154794 696454 155414 706512
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2576 155414 11898
rect 154794 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 155414 -2576
rect 154794 -2896 155414 -2812
rect 154794 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 155414 -2896
rect 154794 -7964 155414 -3132
rect 159294 708028 159914 711900
rect 159294 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 159914 708028
rect 159294 707708 159914 707792
rect 159294 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 159914 707708
rect 159294 700954 159914 707472
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 124954 159914 160398
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3536 159914 16398
rect 159294 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 159914 -3536
rect 159294 -3856 159914 -3772
rect 159294 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 159914 -3856
rect 159294 -7964 159914 -4092
rect 163794 708988 164414 711900
rect 163794 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 164414 708988
rect 163794 708668 164414 708752
rect 163794 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 164414 708668
rect 163794 669454 164414 708432
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4496 164414 20898
rect 163794 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 164414 -4496
rect 163794 -4816 164414 -4732
rect 163794 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 164414 -4816
rect 163794 -7964 164414 -5052
rect 168294 709948 168914 711900
rect 168294 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 168914 709948
rect 168294 709628 168914 709712
rect 168294 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 168914 709628
rect 168294 673954 168914 709392
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5456 168914 25398
rect 168294 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 168914 -5456
rect 168294 -5776 168914 -5692
rect 168294 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 168914 -5776
rect 168294 -7964 168914 -6012
rect 172794 710908 173414 711900
rect 172794 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 173414 710908
rect 172794 710588 173414 710672
rect 172794 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 173414 710588
rect 172794 678454 173414 710352
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6416 173414 29898
rect 172794 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 173414 -6416
rect 172794 -6736 173414 -6652
rect 172794 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 173414 -6736
rect 172794 -7964 173414 -6972
rect 177294 711868 177914 711900
rect 177294 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 177914 711868
rect 177294 711548 177914 711632
rect 177294 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 177914 711548
rect 177294 682954 177914 711312
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7376 177914 34398
rect 177294 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 177914 -7376
rect 177294 -7696 177914 -7612
rect 177294 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 177914 -7696
rect 177294 -7964 177914 -7932
rect 181794 705148 182414 711900
rect 181794 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 182414 705148
rect 181794 704828 182414 704912
rect 181794 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 182414 704828
rect 181794 687454 182414 704592
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -656 182414 2898
rect 181794 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 182414 -656
rect 181794 -976 182414 -892
rect 181794 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 182414 -976
rect 181794 -7964 182414 -1212
rect 186294 706108 186914 711900
rect 186294 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 186914 706108
rect 186294 705788 186914 705872
rect 186294 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 186914 705788
rect 186294 691954 186914 705552
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1616 186914 7398
rect 186294 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 186914 -1616
rect 186294 -1936 186914 -1852
rect 186294 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 186914 -1936
rect 186294 -7964 186914 -2172
rect 190794 707068 191414 711900
rect 190794 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 191414 707068
rect 190794 706748 191414 706832
rect 190794 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 191414 706748
rect 190794 696454 191414 706512
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2576 191414 11898
rect 190794 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 191414 -2576
rect 190794 -2896 191414 -2812
rect 190794 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 191414 -2896
rect 190794 -7964 191414 -3132
rect 195294 708028 195914 711900
rect 195294 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 195914 708028
rect 195294 707708 195914 707792
rect 195294 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 195914 707708
rect 195294 700954 195914 707472
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3536 195914 16398
rect 195294 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 195914 -3536
rect 195294 -3856 195914 -3772
rect 195294 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 195914 -3856
rect 195294 -7964 195914 -4092
rect 199794 708988 200414 711900
rect 199794 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 200414 708988
rect 199794 708668 200414 708752
rect 199794 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 200414 708668
rect 199794 669454 200414 708432
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4496 200414 20898
rect 199794 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 200414 -4496
rect 199794 -4816 200414 -4732
rect 199794 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 200414 -4816
rect 199794 -7964 200414 -5052
rect 204294 709948 204914 711900
rect 204294 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 204914 709948
rect 204294 709628 204914 709712
rect 204294 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 204914 709628
rect 204294 673954 204914 709392
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5456 204914 25398
rect 204294 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 204914 -5456
rect 204294 -5776 204914 -5692
rect 204294 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 204914 -5776
rect 204294 -7964 204914 -6012
rect 208794 710908 209414 711900
rect 208794 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 209414 710908
rect 208794 710588 209414 710672
rect 208794 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 209414 710588
rect 208794 678454 209414 710352
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6416 209414 29898
rect 208794 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 209414 -6416
rect 208794 -6736 209414 -6652
rect 208794 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 209414 -6736
rect 208794 -7964 209414 -6972
rect 213294 711868 213914 711900
rect 213294 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 213914 711868
rect 213294 711548 213914 711632
rect 213294 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 213914 711548
rect 213294 682954 213914 711312
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7376 213914 34398
rect 213294 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 213914 -7376
rect 213294 -7696 213914 -7612
rect 213294 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 213914 -7696
rect 213294 -7964 213914 -7932
rect 217794 705148 218414 711900
rect 217794 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 218414 705148
rect 217794 704828 218414 704912
rect 217794 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 218414 704828
rect 217794 687454 218414 704592
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -656 218414 2898
rect 217794 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 218414 -656
rect 217794 -976 218414 -892
rect 217794 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 218414 -976
rect 217794 -7964 218414 -1212
rect 222294 706108 222914 711900
rect 222294 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 222914 706108
rect 222294 705788 222914 705872
rect 222294 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 222914 705788
rect 222294 691954 222914 705552
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1616 222914 7398
rect 222294 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 222914 -1616
rect 222294 -1936 222914 -1852
rect 222294 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 222914 -1936
rect 222294 -7964 222914 -2172
rect 226794 707068 227414 711900
rect 226794 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 227414 707068
rect 226794 706748 227414 706832
rect 226794 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 227414 706748
rect 226794 696454 227414 706512
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2576 227414 11898
rect 226794 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 227414 -2576
rect 226794 -2896 227414 -2812
rect 226794 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 227414 -2896
rect 226794 -7964 227414 -3132
rect 231294 708028 231914 711900
rect 231294 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 231914 708028
rect 231294 707708 231914 707792
rect 231294 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 231914 707708
rect 231294 700954 231914 707472
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3536 231914 16398
rect 231294 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 231914 -3536
rect 231294 -3856 231914 -3772
rect 231294 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 231914 -3856
rect 231294 -7964 231914 -4092
rect 235794 708988 236414 711900
rect 235794 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 236414 708988
rect 235794 708668 236414 708752
rect 235794 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 236414 708668
rect 235794 669454 236414 708432
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4496 236414 20898
rect 235794 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 236414 -4496
rect 235794 -4816 236414 -4732
rect 235794 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 236414 -4816
rect 235794 -7964 236414 -5052
rect 240294 709948 240914 711900
rect 240294 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 240914 709948
rect 240294 709628 240914 709712
rect 240294 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 240914 709628
rect 240294 673954 240914 709392
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5456 240914 25398
rect 240294 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 240914 -5456
rect 240294 -5776 240914 -5692
rect 240294 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 240914 -5776
rect 240294 -7964 240914 -6012
rect 244794 710908 245414 711900
rect 244794 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 245414 710908
rect 244794 710588 245414 710672
rect 244794 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 245414 710588
rect 244794 678454 245414 710352
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6416 245414 29898
rect 244794 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 245414 -6416
rect 244794 -6736 245414 -6652
rect 244794 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 245414 -6736
rect 244794 -7964 245414 -6972
rect 249294 711868 249914 711900
rect 249294 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 249914 711868
rect 249294 711548 249914 711632
rect 249294 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 249914 711548
rect 249294 682954 249914 711312
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7376 249914 34398
rect 249294 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 249914 -7376
rect 249294 -7696 249914 -7612
rect 249294 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 249914 -7696
rect 249294 -7964 249914 -7932
rect 253794 705148 254414 711900
rect 253794 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 254414 705148
rect 253794 704828 254414 704912
rect 253794 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 254414 704828
rect 253794 687454 254414 704592
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -656 254414 2898
rect 253794 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 254414 -656
rect 253794 -976 254414 -892
rect 253794 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 254414 -976
rect 253794 -7964 254414 -1212
rect 258294 706108 258914 711900
rect 258294 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 258914 706108
rect 258294 705788 258914 705872
rect 258294 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 258914 705788
rect 258294 691954 258914 705552
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1616 258914 7398
rect 258294 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 258914 -1616
rect 258294 -1936 258914 -1852
rect 258294 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 258914 -1936
rect 258294 -7964 258914 -2172
rect 262794 707068 263414 711900
rect 262794 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 263414 707068
rect 262794 706748 263414 706832
rect 262794 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 263414 706748
rect 262794 696454 263414 706512
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2576 263414 11898
rect 262794 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 263414 -2576
rect 262794 -2896 263414 -2812
rect 262794 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 263414 -2896
rect 262794 -7964 263414 -3132
rect 267294 708028 267914 711900
rect 267294 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 267914 708028
rect 267294 707708 267914 707792
rect 267294 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 267914 707708
rect 267294 700954 267914 707472
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3536 267914 16398
rect 267294 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 267914 -3536
rect 267294 -3856 267914 -3772
rect 267294 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 267914 -3856
rect 267294 -7964 267914 -4092
rect 271794 708988 272414 711900
rect 271794 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 272414 708988
rect 271794 708668 272414 708752
rect 271794 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 272414 708668
rect 271794 669454 272414 708432
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4496 272414 20898
rect 271794 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 272414 -4496
rect 271794 -4816 272414 -4732
rect 271794 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 272414 -4816
rect 271794 -7964 272414 -5052
rect 276294 709948 276914 711900
rect 276294 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 276914 709948
rect 276294 709628 276914 709712
rect 276294 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 276914 709628
rect 276294 673954 276914 709392
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5456 276914 25398
rect 276294 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 276914 -5456
rect 276294 -5776 276914 -5692
rect 276294 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 276914 -5776
rect 276294 -7964 276914 -6012
rect 280794 710908 281414 711900
rect 280794 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 281414 710908
rect 280794 710588 281414 710672
rect 280794 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 281414 710588
rect 280794 678454 281414 710352
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6416 281414 29898
rect 280794 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 281414 -6416
rect 280794 -6736 281414 -6652
rect 280794 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 281414 -6736
rect 280794 -7964 281414 -6972
rect 285294 711868 285914 711900
rect 285294 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 285914 711868
rect 285294 711548 285914 711632
rect 285294 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 285914 711548
rect 285294 682954 285914 711312
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7376 285914 34398
rect 285294 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 285914 -7376
rect 285294 -7696 285914 -7612
rect 285294 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 285914 -7696
rect 285294 -7964 285914 -7932
rect 289794 705148 290414 711900
rect 289794 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 290414 705148
rect 289794 704828 290414 704912
rect 289794 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 290414 704828
rect 289794 687454 290414 704592
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -656 290414 2898
rect 289794 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 290414 -656
rect 289794 -976 290414 -892
rect 289794 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 290414 -976
rect 289794 -7964 290414 -1212
rect 294294 706108 294914 711900
rect 294294 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 294914 706108
rect 294294 705788 294914 705872
rect 294294 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 294914 705788
rect 294294 691954 294914 705552
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1616 294914 7398
rect 294294 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 294914 -1616
rect 294294 -1936 294914 -1852
rect 294294 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 294914 -1936
rect 294294 -7964 294914 -2172
rect 298794 707068 299414 711900
rect 298794 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 299414 707068
rect 298794 706748 299414 706832
rect 298794 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 299414 706748
rect 298794 696454 299414 706512
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2576 299414 11898
rect 298794 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 299414 -2576
rect 298794 -2896 299414 -2812
rect 298794 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 299414 -2896
rect 298794 -7964 299414 -3132
rect 303294 708028 303914 711900
rect 303294 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 303914 708028
rect 303294 707708 303914 707792
rect 303294 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 303914 707708
rect 303294 700954 303914 707472
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3536 303914 16398
rect 303294 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 303914 -3536
rect 303294 -3856 303914 -3772
rect 303294 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 303914 -3856
rect 303294 -7964 303914 -4092
rect 307794 708988 308414 711900
rect 307794 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 308414 708988
rect 307794 708668 308414 708752
rect 307794 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 308414 708668
rect 307794 669454 308414 708432
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4496 308414 20898
rect 307794 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 308414 -4496
rect 307794 -4816 308414 -4732
rect 307794 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 308414 -4816
rect 307794 -7964 308414 -5052
rect 312294 709948 312914 711900
rect 312294 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 312914 709948
rect 312294 709628 312914 709712
rect 312294 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 312914 709628
rect 312294 673954 312914 709392
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5456 312914 25398
rect 312294 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 312914 -5456
rect 312294 -5776 312914 -5692
rect 312294 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 312914 -5776
rect 312294 -7964 312914 -6012
rect 316794 710908 317414 711900
rect 316794 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 317414 710908
rect 316794 710588 317414 710672
rect 316794 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 317414 710588
rect 316794 678454 317414 710352
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6416 317414 29898
rect 316794 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 317414 -6416
rect 316794 -6736 317414 -6652
rect 316794 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 317414 -6736
rect 316794 -7964 317414 -6972
rect 321294 711868 321914 711900
rect 321294 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 321914 711868
rect 321294 711548 321914 711632
rect 321294 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 321914 711548
rect 321294 682954 321914 711312
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7376 321914 34398
rect 321294 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 321914 -7376
rect 321294 -7696 321914 -7612
rect 321294 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 321914 -7696
rect 321294 -7964 321914 -7932
rect 325794 705148 326414 711900
rect 325794 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 326414 705148
rect 325794 704828 326414 704912
rect 325794 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 326414 704828
rect 325794 687454 326414 704592
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -656 326414 2898
rect 325794 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 326414 -656
rect 325794 -976 326414 -892
rect 325794 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 326414 -976
rect 325794 -7964 326414 -1212
rect 330294 706108 330914 711900
rect 330294 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 330914 706108
rect 330294 705788 330914 705872
rect 330294 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 330914 705788
rect 330294 691954 330914 705552
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1616 330914 7398
rect 330294 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 330914 -1616
rect 330294 -1936 330914 -1852
rect 330294 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 330914 -1936
rect 330294 -7964 330914 -2172
rect 334794 707068 335414 711900
rect 334794 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 335414 707068
rect 334794 706748 335414 706832
rect 334794 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 335414 706748
rect 334794 696454 335414 706512
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2576 335414 11898
rect 334794 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 335414 -2576
rect 334794 -2896 335414 -2812
rect 334794 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 335414 -2896
rect 334794 -7964 335414 -3132
rect 339294 708028 339914 711900
rect 339294 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 339914 708028
rect 339294 707708 339914 707792
rect 339294 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 339914 707708
rect 339294 700954 339914 707472
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3536 339914 16398
rect 339294 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 339914 -3536
rect 339294 -3856 339914 -3772
rect 339294 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 339914 -3856
rect 339294 -7964 339914 -4092
rect 343794 708988 344414 711900
rect 343794 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 344414 708988
rect 343794 708668 344414 708752
rect 343794 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 344414 708668
rect 343794 669454 344414 708432
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4496 344414 20898
rect 343794 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 344414 -4496
rect 343794 -4816 344414 -4732
rect 343794 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 344414 -4816
rect 343794 -7964 344414 -5052
rect 348294 709948 348914 711900
rect 348294 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 348914 709948
rect 348294 709628 348914 709712
rect 348294 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 348914 709628
rect 348294 673954 348914 709392
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5456 348914 25398
rect 348294 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 348914 -5456
rect 348294 -5776 348914 -5692
rect 348294 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 348914 -5776
rect 348294 -7964 348914 -6012
rect 352794 710908 353414 711900
rect 352794 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 353414 710908
rect 352794 710588 353414 710672
rect 352794 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 353414 710588
rect 352794 678454 353414 710352
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6416 353414 29898
rect 352794 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 353414 -6416
rect 352794 -6736 353414 -6652
rect 352794 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 353414 -6736
rect 352794 -7964 353414 -6972
rect 357294 711868 357914 711900
rect 357294 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 357914 711868
rect 357294 711548 357914 711632
rect 357294 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 357914 711548
rect 357294 682954 357914 711312
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7376 357914 34398
rect 357294 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 357914 -7376
rect 357294 -7696 357914 -7612
rect 357294 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 357914 -7696
rect 357294 -7964 357914 -7932
rect 361794 705148 362414 711900
rect 361794 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 362414 705148
rect 361794 704828 362414 704912
rect 361794 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 362414 704828
rect 361794 687454 362414 704592
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -656 362414 2898
rect 361794 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 362414 -656
rect 361794 -976 362414 -892
rect 361794 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 362414 -976
rect 361794 -7964 362414 -1212
rect 366294 706108 366914 711900
rect 366294 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 366914 706108
rect 366294 705788 366914 705872
rect 366294 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 366914 705788
rect 366294 691954 366914 705552
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1616 366914 7398
rect 366294 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 366914 -1616
rect 366294 -1936 366914 -1852
rect 366294 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 366914 -1936
rect 366294 -7964 366914 -2172
rect 370794 707068 371414 711900
rect 370794 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 371414 707068
rect 370794 706748 371414 706832
rect 370794 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 371414 706748
rect 370794 696454 371414 706512
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2576 371414 11898
rect 370794 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 371414 -2576
rect 370794 -2896 371414 -2812
rect 370794 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 371414 -2896
rect 370794 -7964 371414 -3132
rect 375294 708028 375914 711900
rect 375294 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 375914 708028
rect 375294 707708 375914 707792
rect 375294 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 375914 707708
rect 375294 700954 375914 707472
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3536 375914 16398
rect 375294 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 375914 -3536
rect 375294 -3856 375914 -3772
rect 375294 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 375914 -3856
rect 375294 -7964 375914 -4092
rect 379794 708988 380414 711900
rect 379794 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 380414 708988
rect 379794 708668 380414 708752
rect 379794 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 380414 708668
rect 379794 669454 380414 708432
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4496 380414 20898
rect 379794 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 380414 -4496
rect 379794 -4816 380414 -4732
rect 379794 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 380414 -4816
rect 379794 -7964 380414 -5052
rect 384294 709948 384914 711900
rect 384294 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 384914 709948
rect 384294 709628 384914 709712
rect 384294 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 384914 709628
rect 384294 673954 384914 709392
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5456 384914 25398
rect 384294 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 384914 -5456
rect 384294 -5776 384914 -5692
rect 384294 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 384914 -5776
rect 384294 -7964 384914 -6012
rect 388794 710908 389414 711900
rect 388794 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 389414 710908
rect 388794 710588 389414 710672
rect 388794 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 389414 710588
rect 388794 678454 389414 710352
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6416 389414 29898
rect 388794 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 389414 -6416
rect 388794 -6736 389414 -6652
rect 388794 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 389414 -6736
rect 388794 -7964 389414 -6972
rect 393294 711868 393914 711900
rect 393294 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 393914 711868
rect 393294 711548 393914 711632
rect 393294 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 393914 711548
rect 393294 682954 393914 711312
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7376 393914 34398
rect 393294 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 393914 -7376
rect 393294 -7696 393914 -7612
rect 393294 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 393914 -7696
rect 393294 -7964 393914 -7932
rect 397794 705148 398414 711900
rect 397794 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 398414 705148
rect 397794 704828 398414 704912
rect 397794 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 398414 704828
rect 397794 687454 398414 704592
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -656 398414 2898
rect 397794 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 398414 -656
rect 397794 -976 398414 -892
rect 397794 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 398414 -976
rect 397794 -7964 398414 -1212
rect 402294 706108 402914 711900
rect 402294 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 402914 706108
rect 402294 705788 402914 705872
rect 402294 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 402914 705788
rect 402294 691954 402914 705552
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1616 402914 7398
rect 402294 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 402914 -1616
rect 402294 -1936 402914 -1852
rect 402294 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 402914 -1936
rect 402294 -7964 402914 -2172
rect 406794 707068 407414 711900
rect 406794 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 407414 707068
rect 406794 706748 407414 706832
rect 406794 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 407414 706748
rect 406794 696454 407414 706512
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2576 407414 11898
rect 406794 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 407414 -2576
rect 406794 -2896 407414 -2812
rect 406794 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 407414 -2896
rect 406794 -7964 407414 -3132
rect 411294 708028 411914 711900
rect 411294 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 411914 708028
rect 411294 707708 411914 707792
rect 411294 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 411914 707708
rect 411294 700954 411914 707472
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3536 411914 16398
rect 411294 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 411914 -3536
rect 411294 -3856 411914 -3772
rect 411294 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 411914 -3856
rect 411294 -7964 411914 -4092
rect 415794 708988 416414 711900
rect 415794 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 416414 708988
rect 415794 708668 416414 708752
rect 415794 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 416414 708668
rect 415794 669454 416414 708432
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4496 416414 20898
rect 415794 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 416414 -4496
rect 415794 -4816 416414 -4732
rect 415794 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 416414 -4816
rect 415794 -7964 416414 -5052
rect 420294 709948 420914 711900
rect 420294 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 420914 709948
rect 420294 709628 420914 709712
rect 420294 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 420914 709628
rect 420294 673954 420914 709392
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5456 420914 25398
rect 420294 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 420914 -5456
rect 420294 -5776 420914 -5692
rect 420294 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 420914 -5776
rect 420294 -7964 420914 -6012
rect 424794 710908 425414 711900
rect 424794 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 425414 710908
rect 424794 710588 425414 710672
rect 424794 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 425414 710588
rect 424794 678454 425414 710352
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6416 425414 29898
rect 424794 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 425414 -6416
rect 424794 -6736 425414 -6652
rect 424794 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 425414 -6736
rect 424794 -7964 425414 -6972
rect 429294 711868 429914 711900
rect 429294 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 429914 711868
rect 429294 711548 429914 711632
rect 429294 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 429914 711548
rect 429294 682954 429914 711312
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7376 429914 34398
rect 429294 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 429914 -7376
rect 429294 -7696 429914 -7612
rect 429294 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 429914 -7696
rect 429294 -7964 429914 -7932
rect 433794 705148 434414 711900
rect 433794 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 434414 705148
rect 433794 704828 434414 704912
rect 433794 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 434414 704828
rect 433794 687454 434414 704592
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -656 434414 2898
rect 433794 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 434414 -656
rect 433794 -976 434414 -892
rect 433794 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 434414 -976
rect 433794 -7964 434414 -1212
rect 438294 706108 438914 711900
rect 438294 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 438914 706108
rect 438294 705788 438914 705872
rect 438294 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 438914 705788
rect 438294 691954 438914 705552
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1616 438914 7398
rect 438294 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 438914 -1616
rect 438294 -1936 438914 -1852
rect 438294 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 438914 -1936
rect 438294 -7964 438914 -2172
rect 442794 707068 443414 711900
rect 442794 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 443414 707068
rect 442794 706748 443414 706832
rect 442794 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 443414 706748
rect 442794 696454 443414 706512
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2576 443414 11898
rect 442794 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 443414 -2576
rect 442794 -2896 443414 -2812
rect 442794 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 443414 -2896
rect 442794 -7964 443414 -3132
rect 447294 708028 447914 711900
rect 447294 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 447914 708028
rect 447294 707708 447914 707792
rect 447294 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 447914 707708
rect 447294 700954 447914 707472
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3536 447914 16398
rect 447294 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 447914 -3536
rect 447294 -3856 447914 -3772
rect 447294 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 447914 -3856
rect 447294 -7964 447914 -4092
rect 451794 708988 452414 711900
rect 451794 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 452414 708988
rect 451794 708668 452414 708752
rect 451794 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 452414 708668
rect 451794 669454 452414 708432
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4496 452414 20898
rect 451794 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 452414 -4496
rect 451794 -4816 452414 -4732
rect 451794 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 452414 -4816
rect 451794 -7964 452414 -5052
rect 456294 709948 456914 711900
rect 456294 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 456914 709948
rect 456294 709628 456914 709712
rect 456294 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 456914 709628
rect 456294 673954 456914 709392
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5456 456914 25398
rect 456294 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 456914 -5456
rect 456294 -5776 456914 -5692
rect 456294 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 456914 -5776
rect 456294 -7964 456914 -6012
rect 460794 710908 461414 711900
rect 460794 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 461414 710908
rect 460794 710588 461414 710672
rect 460794 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 461414 710588
rect 460794 678454 461414 710352
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6416 461414 29898
rect 460794 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 461414 -6416
rect 460794 -6736 461414 -6652
rect 460794 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 461414 -6736
rect 460794 -7964 461414 -6972
rect 465294 711868 465914 711900
rect 465294 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 465914 711868
rect 465294 711548 465914 711632
rect 465294 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 465914 711548
rect 465294 682954 465914 711312
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7376 465914 34398
rect 465294 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 465914 -7376
rect 465294 -7696 465914 -7612
rect 465294 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 465914 -7696
rect 465294 -7964 465914 -7932
rect 469794 705148 470414 711900
rect 469794 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 470414 705148
rect 469794 704828 470414 704912
rect 469794 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 470414 704828
rect 469794 687454 470414 704592
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -656 470414 2898
rect 469794 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 470414 -656
rect 469794 -976 470414 -892
rect 469794 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 470414 -976
rect 469794 -7964 470414 -1212
rect 474294 706108 474914 711900
rect 474294 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 474914 706108
rect 474294 705788 474914 705872
rect 474294 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 474914 705788
rect 474294 691954 474914 705552
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1616 474914 7398
rect 474294 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 474914 -1616
rect 474294 -1936 474914 -1852
rect 474294 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 474914 -1936
rect 474294 -7964 474914 -2172
rect 478794 707068 479414 711900
rect 478794 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 479414 707068
rect 478794 706748 479414 706832
rect 478794 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 479414 706748
rect 478794 696454 479414 706512
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2576 479414 11898
rect 478794 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 479414 -2576
rect 478794 -2896 479414 -2812
rect 478794 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 479414 -2896
rect 478794 -7964 479414 -3132
rect 483294 708028 483914 711900
rect 483294 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 483914 708028
rect 483294 707708 483914 707792
rect 483294 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 483914 707708
rect 483294 700954 483914 707472
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3536 483914 16398
rect 483294 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 483914 -3536
rect 483294 -3856 483914 -3772
rect 483294 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 483914 -3856
rect 483294 -7964 483914 -4092
rect 487794 708988 488414 711900
rect 487794 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 488414 708988
rect 487794 708668 488414 708752
rect 487794 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 488414 708668
rect 487794 669454 488414 708432
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4496 488414 20898
rect 487794 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 488414 -4496
rect 487794 -4816 488414 -4732
rect 487794 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 488414 -4816
rect 487794 -7964 488414 -5052
rect 492294 709948 492914 711900
rect 492294 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 492914 709948
rect 492294 709628 492914 709712
rect 492294 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 492914 709628
rect 492294 673954 492914 709392
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5456 492914 25398
rect 492294 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 492914 -5456
rect 492294 -5776 492914 -5692
rect 492294 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 492914 -5776
rect 492294 -7964 492914 -6012
rect 496794 710908 497414 711900
rect 496794 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 497414 710908
rect 496794 710588 497414 710672
rect 496794 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 497414 710588
rect 496794 678454 497414 710352
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6416 497414 29898
rect 496794 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 497414 -6416
rect 496794 -6736 497414 -6652
rect 496794 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 497414 -6736
rect 496794 -7964 497414 -6972
rect 501294 711868 501914 711900
rect 501294 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 501914 711868
rect 501294 711548 501914 711632
rect 501294 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 501914 711548
rect 501294 682954 501914 711312
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7376 501914 34398
rect 501294 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 501914 -7376
rect 501294 -7696 501914 -7612
rect 501294 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 501914 -7696
rect 501294 -7964 501914 -7932
rect 505794 705148 506414 711900
rect 505794 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 506414 705148
rect 505794 704828 506414 704912
rect 505794 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 506414 704828
rect 505794 687454 506414 704592
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -656 506414 2898
rect 505794 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 506414 -656
rect 505794 -976 506414 -892
rect 505794 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 506414 -976
rect 505794 -7964 506414 -1212
rect 510294 706108 510914 711900
rect 510294 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 510914 706108
rect 510294 705788 510914 705872
rect 510294 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 510914 705788
rect 510294 691954 510914 705552
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1616 510914 7398
rect 510294 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 510914 -1616
rect 510294 -1936 510914 -1852
rect 510294 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 510914 -1936
rect 510294 -7964 510914 -2172
rect 514794 707068 515414 711900
rect 514794 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 515414 707068
rect 514794 706748 515414 706832
rect 514794 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 515414 706748
rect 514794 696454 515414 706512
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2576 515414 11898
rect 514794 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 515414 -2576
rect 514794 -2896 515414 -2812
rect 514794 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 515414 -2896
rect 514794 -7964 515414 -3132
rect 519294 708028 519914 711900
rect 519294 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 519914 708028
rect 519294 707708 519914 707792
rect 519294 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 519914 707708
rect 519294 700954 519914 707472
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3536 519914 16398
rect 519294 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 519914 -3536
rect 519294 -3856 519914 -3772
rect 519294 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 519914 -3856
rect 519294 -7964 519914 -4092
rect 523794 708988 524414 711900
rect 523794 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 524414 708988
rect 523794 708668 524414 708752
rect 523794 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 524414 708668
rect 523794 669454 524414 708432
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4496 524414 20898
rect 523794 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 524414 -4496
rect 523794 -4816 524414 -4732
rect 523794 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 524414 -4816
rect 523794 -7964 524414 -5052
rect 528294 709948 528914 711900
rect 528294 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 528914 709948
rect 528294 709628 528914 709712
rect 528294 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 528914 709628
rect 528294 673954 528914 709392
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5456 528914 25398
rect 528294 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 528914 -5456
rect 528294 -5776 528914 -5692
rect 528294 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 528914 -5776
rect 528294 -7964 528914 -6012
rect 532794 710908 533414 711900
rect 532794 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 533414 710908
rect 532794 710588 533414 710672
rect 532794 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 533414 710588
rect 532794 678454 533414 710352
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6416 533414 29898
rect 532794 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 533414 -6416
rect 532794 -6736 533414 -6652
rect 532794 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 533414 -6736
rect 532794 -7964 533414 -6972
rect 537294 711868 537914 711900
rect 537294 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 537914 711868
rect 537294 711548 537914 711632
rect 537294 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 537914 711548
rect 537294 682954 537914 711312
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7376 537914 34398
rect 537294 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 537914 -7376
rect 537294 -7696 537914 -7612
rect 537294 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 537914 -7696
rect 537294 -7964 537914 -7932
rect 541794 705148 542414 711900
rect 541794 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 542414 705148
rect 541794 704828 542414 704912
rect 541794 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 542414 704828
rect 541794 687454 542414 704592
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -656 542414 2898
rect 541794 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 542414 -656
rect 541794 -976 542414 -892
rect 541794 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 542414 -976
rect 541794 -7964 542414 -1212
rect 546294 706108 546914 711900
rect 546294 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 546914 706108
rect 546294 705788 546914 705872
rect 546294 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 546914 705788
rect 546294 691954 546914 705552
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1616 546914 7398
rect 546294 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 546914 -1616
rect 546294 -1936 546914 -1852
rect 546294 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 546914 -1936
rect 546294 -7964 546914 -2172
rect 550794 707068 551414 711900
rect 550794 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 551414 707068
rect 550794 706748 551414 706832
rect 550794 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 551414 706748
rect 550794 696454 551414 706512
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2576 551414 11898
rect 550794 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 551414 -2576
rect 550794 -2896 551414 -2812
rect 550794 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 551414 -2896
rect 550794 -7964 551414 -3132
rect 555294 708028 555914 711900
rect 555294 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 555914 708028
rect 555294 707708 555914 707792
rect 555294 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 555914 707708
rect 555294 700954 555914 707472
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3536 555914 16398
rect 555294 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 555914 -3536
rect 555294 -3856 555914 -3772
rect 555294 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 555914 -3856
rect 555294 -7964 555914 -4092
rect 559794 708988 560414 711900
rect 559794 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 560414 708988
rect 559794 708668 560414 708752
rect 559794 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 560414 708668
rect 559794 669454 560414 708432
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4496 560414 20898
rect 559794 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 560414 -4496
rect 559794 -4816 560414 -4732
rect 559794 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 560414 -4816
rect 559794 -7964 560414 -5052
rect 564294 709948 564914 711900
rect 564294 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 564914 709948
rect 564294 709628 564914 709712
rect 564294 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 564914 709628
rect 564294 673954 564914 709392
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5456 564914 25398
rect 564294 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 564914 -5456
rect 564294 -5776 564914 -5692
rect 564294 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 564914 -5776
rect 564294 -7964 564914 -6012
rect 568794 710908 569414 711900
rect 568794 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 569414 710908
rect 568794 710588 569414 710672
rect 568794 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 569414 710588
rect 568794 678454 569414 710352
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6416 569414 29898
rect 568794 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 569414 -6416
rect 568794 -6736 569414 -6652
rect 568794 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 569414 -6736
rect 568794 -7964 569414 -6972
rect 573294 711868 573914 711900
rect 573294 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 573914 711868
rect 573294 711548 573914 711632
rect 573294 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 573914 711548
rect 573294 682954 573914 711312
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7376 573914 34398
rect 573294 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 573914 -7376
rect 573294 -7696 573914 -7612
rect 573294 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 573914 -7696
rect 573294 -7964 573914 -7932
rect 577794 705148 578414 711900
rect 577794 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 578414 705148
rect 577794 704828 578414 704912
rect 577794 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 578414 704828
rect 577794 687454 578414 704592
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -656 578414 2898
rect 577794 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 578414 -656
rect 577794 -976 578414 -892
rect 577794 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 578414 -976
rect 577794 -7964 578414 -1212
rect 582294 706108 582914 711900
rect 592340 711868 592960 711900
rect 592340 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect 592340 711548 592960 711632
rect 592340 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect 591380 710908 592000 710940
rect 591380 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect 591380 710588 592000 710672
rect 591380 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect 590420 709948 591040 709980
rect 590420 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect 590420 709628 591040 709712
rect 590420 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect 589460 708988 590080 709020
rect 589460 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect 589460 708668 590080 708752
rect 589460 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect 588500 708028 589120 708060
rect 588500 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect 588500 707708 589120 707792
rect 588500 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect 587540 707068 588160 707100
rect 587540 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect 587540 706748 588160 706832
rect 587540 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect 582294 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 582914 706108
rect 582294 705788 582914 705872
rect 582294 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 582914 705788
rect 582294 691954 582914 705552
rect 586580 706108 587200 706140
rect 586580 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect 586580 705788 587200 705872
rect 586580 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1616 582914 7398
rect 585620 705148 586240 705180
rect 585620 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect 585620 704828 586240 704912
rect 585620 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect 585620 687454 586240 704592
rect 585620 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 586240 687454
rect 585620 687134 586240 687218
rect 585620 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 586240 687134
rect 585620 651454 586240 686898
rect 585620 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 586240 651454
rect 585620 651134 586240 651218
rect 585620 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 586240 651134
rect 585620 615454 586240 650898
rect 585620 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 586240 615454
rect 585620 615134 586240 615218
rect 585620 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 586240 615134
rect 585620 579454 586240 614898
rect 585620 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 586240 579454
rect 585620 579134 586240 579218
rect 585620 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 586240 579134
rect 585620 543454 586240 578898
rect 585620 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 586240 543454
rect 585620 543134 586240 543218
rect 585620 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 586240 543134
rect 585620 507454 586240 542898
rect 585620 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 586240 507454
rect 585620 507134 586240 507218
rect 585620 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 586240 507134
rect 585620 471454 586240 506898
rect 585620 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 586240 471454
rect 585620 471134 586240 471218
rect 585620 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 586240 471134
rect 585620 435454 586240 470898
rect 585620 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 586240 435454
rect 585620 435134 586240 435218
rect 585620 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 586240 435134
rect 585620 399454 586240 434898
rect 585620 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 586240 399454
rect 585620 399134 586240 399218
rect 585620 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 586240 399134
rect 585620 363454 586240 398898
rect 585620 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 586240 363454
rect 585620 363134 586240 363218
rect 585620 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 586240 363134
rect 585620 327454 586240 362898
rect 585620 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 586240 327454
rect 585620 327134 586240 327218
rect 585620 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 586240 327134
rect 585620 291454 586240 326898
rect 585620 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 586240 291454
rect 585620 291134 586240 291218
rect 585620 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 586240 291134
rect 585620 255454 586240 290898
rect 585620 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 586240 255454
rect 585620 255134 586240 255218
rect 585620 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 586240 255134
rect 585620 219454 586240 254898
rect 585620 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 586240 219454
rect 585620 219134 586240 219218
rect 585620 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 586240 219134
rect 585620 183454 586240 218898
rect 585620 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 586240 183454
rect 585620 183134 586240 183218
rect 585620 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 586240 183134
rect 585620 147454 586240 182898
rect 585620 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 586240 147454
rect 585620 147134 586240 147218
rect 585620 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 586240 147134
rect 585620 111454 586240 146898
rect 585620 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 586240 111454
rect 585620 111134 586240 111218
rect 585620 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 586240 111134
rect 585620 75454 586240 110898
rect 585620 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 586240 75454
rect 585620 75134 586240 75218
rect 585620 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 586240 75134
rect 585620 39454 586240 74898
rect 585620 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 586240 39454
rect 585620 39134 586240 39218
rect 585620 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 586240 39134
rect 585620 3454 586240 38898
rect 585620 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 586240 3454
rect 585620 3134 586240 3218
rect 585620 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 586240 3134
rect 585620 -656 586240 2898
rect 585620 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect 585620 -976 586240 -892
rect 585620 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect 585620 -1244 586240 -1212
rect 586580 691954 587200 705552
rect 586580 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 587200 691954
rect 586580 691634 587200 691718
rect 586580 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 587200 691634
rect 586580 655954 587200 691398
rect 586580 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 587200 655954
rect 586580 655634 587200 655718
rect 586580 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 587200 655634
rect 586580 619954 587200 655398
rect 586580 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 587200 619954
rect 586580 619634 587200 619718
rect 586580 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 587200 619634
rect 586580 583954 587200 619398
rect 586580 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 587200 583954
rect 586580 583634 587200 583718
rect 586580 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 587200 583634
rect 586580 547954 587200 583398
rect 586580 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 587200 547954
rect 586580 547634 587200 547718
rect 586580 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 587200 547634
rect 586580 511954 587200 547398
rect 586580 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 587200 511954
rect 586580 511634 587200 511718
rect 586580 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 587200 511634
rect 586580 475954 587200 511398
rect 586580 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 587200 475954
rect 586580 475634 587200 475718
rect 586580 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 587200 475634
rect 586580 439954 587200 475398
rect 586580 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 587200 439954
rect 586580 439634 587200 439718
rect 586580 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 587200 439634
rect 586580 403954 587200 439398
rect 586580 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 587200 403954
rect 586580 403634 587200 403718
rect 586580 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 587200 403634
rect 586580 367954 587200 403398
rect 586580 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 587200 367954
rect 586580 367634 587200 367718
rect 586580 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 587200 367634
rect 586580 331954 587200 367398
rect 586580 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 587200 331954
rect 586580 331634 587200 331718
rect 586580 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 587200 331634
rect 586580 295954 587200 331398
rect 586580 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 587200 295954
rect 586580 295634 587200 295718
rect 586580 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 587200 295634
rect 586580 259954 587200 295398
rect 586580 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 587200 259954
rect 586580 259634 587200 259718
rect 586580 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 587200 259634
rect 586580 223954 587200 259398
rect 586580 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 587200 223954
rect 586580 223634 587200 223718
rect 586580 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 587200 223634
rect 586580 187954 587200 223398
rect 586580 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 587200 187954
rect 586580 187634 587200 187718
rect 586580 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 587200 187634
rect 586580 151954 587200 187398
rect 586580 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 587200 151954
rect 586580 151634 587200 151718
rect 586580 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 587200 151634
rect 586580 115954 587200 151398
rect 586580 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 587200 115954
rect 586580 115634 587200 115718
rect 586580 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 587200 115634
rect 586580 79954 587200 115398
rect 586580 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 587200 79954
rect 586580 79634 587200 79718
rect 586580 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 587200 79634
rect 586580 43954 587200 79398
rect 586580 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 587200 43954
rect 586580 43634 587200 43718
rect 586580 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 587200 43634
rect 586580 7954 587200 43398
rect 586580 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 587200 7954
rect 586580 7634 587200 7718
rect 586580 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 587200 7634
rect 582294 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 582914 -1616
rect 582294 -1936 582914 -1852
rect 582294 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 582914 -1936
rect 582294 -7964 582914 -2172
rect 586580 -1616 587200 7398
rect 586580 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect 586580 -1936 587200 -1852
rect 586580 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect 586580 -2204 587200 -2172
rect 587540 696454 588160 706512
rect 587540 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 588160 696454
rect 587540 696134 588160 696218
rect 587540 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 588160 696134
rect 587540 660454 588160 695898
rect 587540 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 588160 660454
rect 587540 660134 588160 660218
rect 587540 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 588160 660134
rect 587540 624454 588160 659898
rect 587540 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 588160 624454
rect 587540 624134 588160 624218
rect 587540 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 588160 624134
rect 587540 588454 588160 623898
rect 587540 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 588160 588454
rect 587540 588134 588160 588218
rect 587540 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 588160 588134
rect 587540 552454 588160 587898
rect 587540 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 588160 552454
rect 587540 552134 588160 552218
rect 587540 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 588160 552134
rect 587540 516454 588160 551898
rect 587540 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 588160 516454
rect 587540 516134 588160 516218
rect 587540 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 588160 516134
rect 587540 480454 588160 515898
rect 587540 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 588160 480454
rect 587540 480134 588160 480218
rect 587540 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 588160 480134
rect 587540 444454 588160 479898
rect 587540 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 588160 444454
rect 587540 444134 588160 444218
rect 587540 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 588160 444134
rect 587540 408454 588160 443898
rect 587540 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 588160 408454
rect 587540 408134 588160 408218
rect 587540 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 588160 408134
rect 587540 372454 588160 407898
rect 587540 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 588160 372454
rect 587540 372134 588160 372218
rect 587540 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 588160 372134
rect 587540 336454 588160 371898
rect 587540 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 588160 336454
rect 587540 336134 588160 336218
rect 587540 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 588160 336134
rect 587540 300454 588160 335898
rect 587540 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 588160 300454
rect 587540 300134 588160 300218
rect 587540 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 588160 300134
rect 587540 264454 588160 299898
rect 587540 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 588160 264454
rect 587540 264134 588160 264218
rect 587540 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 588160 264134
rect 587540 228454 588160 263898
rect 587540 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 588160 228454
rect 587540 228134 588160 228218
rect 587540 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 588160 228134
rect 587540 192454 588160 227898
rect 587540 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 588160 192454
rect 587540 192134 588160 192218
rect 587540 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 588160 192134
rect 587540 156454 588160 191898
rect 587540 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 588160 156454
rect 587540 156134 588160 156218
rect 587540 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 588160 156134
rect 587540 120454 588160 155898
rect 587540 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 588160 120454
rect 587540 120134 588160 120218
rect 587540 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 588160 120134
rect 587540 84454 588160 119898
rect 587540 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 588160 84454
rect 587540 84134 588160 84218
rect 587540 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 588160 84134
rect 587540 48454 588160 83898
rect 587540 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 588160 48454
rect 587540 48134 588160 48218
rect 587540 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 588160 48134
rect 587540 12454 588160 47898
rect 587540 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 588160 12454
rect 587540 12134 588160 12218
rect 587540 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 588160 12134
rect 587540 -2576 588160 11898
rect 587540 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect 587540 -2896 588160 -2812
rect 587540 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect 587540 -3164 588160 -3132
rect 588500 700954 589120 707472
rect 588500 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 589120 700954
rect 588500 700634 589120 700718
rect 588500 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 589120 700634
rect 588500 664954 589120 700398
rect 588500 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 589120 664954
rect 588500 664634 589120 664718
rect 588500 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 589120 664634
rect 588500 628954 589120 664398
rect 588500 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 589120 628954
rect 588500 628634 589120 628718
rect 588500 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 589120 628634
rect 588500 592954 589120 628398
rect 588500 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 589120 592954
rect 588500 592634 589120 592718
rect 588500 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 589120 592634
rect 588500 556954 589120 592398
rect 588500 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 589120 556954
rect 588500 556634 589120 556718
rect 588500 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 589120 556634
rect 588500 520954 589120 556398
rect 588500 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 589120 520954
rect 588500 520634 589120 520718
rect 588500 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 589120 520634
rect 588500 484954 589120 520398
rect 588500 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 589120 484954
rect 588500 484634 589120 484718
rect 588500 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 589120 484634
rect 588500 448954 589120 484398
rect 588500 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 589120 448954
rect 588500 448634 589120 448718
rect 588500 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 589120 448634
rect 588500 412954 589120 448398
rect 588500 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 589120 412954
rect 588500 412634 589120 412718
rect 588500 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 589120 412634
rect 588500 376954 589120 412398
rect 588500 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 589120 376954
rect 588500 376634 589120 376718
rect 588500 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 589120 376634
rect 588500 340954 589120 376398
rect 588500 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 589120 340954
rect 588500 340634 589120 340718
rect 588500 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 589120 340634
rect 588500 304954 589120 340398
rect 588500 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 589120 304954
rect 588500 304634 589120 304718
rect 588500 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 589120 304634
rect 588500 268954 589120 304398
rect 588500 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 589120 268954
rect 588500 268634 589120 268718
rect 588500 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 589120 268634
rect 588500 232954 589120 268398
rect 588500 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 589120 232954
rect 588500 232634 589120 232718
rect 588500 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 589120 232634
rect 588500 196954 589120 232398
rect 588500 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 589120 196954
rect 588500 196634 589120 196718
rect 588500 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 589120 196634
rect 588500 160954 589120 196398
rect 588500 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 589120 160954
rect 588500 160634 589120 160718
rect 588500 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 589120 160634
rect 588500 124954 589120 160398
rect 588500 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 589120 124954
rect 588500 124634 589120 124718
rect 588500 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 589120 124634
rect 588500 88954 589120 124398
rect 588500 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 589120 88954
rect 588500 88634 589120 88718
rect 588500 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 589120 88634
rect 588500 52954 589120 88398
rect 588500 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 589120 52954
rect 588500 52634 589120 52718
rect 588500 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 589120 52634
rect 588500 16954 589120 52398
rect 588500 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 589120 16954
rect 588500 16634 589120 16718
rect 588500 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 589120 16634
rect 588500 -3536 589120 16398
rect 588500 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect 588500 -3856 589120 -3772
rect 588500 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect 588500 -4124 589120 -4092
rect 589460 669454 590080 708432
rect 589460 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 590080 669454
rect 589460 669134 590080 669218
rect 589460 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 590080 669134
rect 589460 633454 590080 668898
rect 589460 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 590080 633454
rect 589460 633134 590080 633218
rect 589460 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 590080 633134
rect 589460 597454 590080 632898
rect 589460 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 590080 597454
rect 589460 597134 590080 597218
rect 589460 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 590080 597134
rect 589460 561454 590080 596898
rect 589460 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 590080 561454
rect 589460 561134 590080 561218
rect 589460 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 590080 561134
rect 589460 525454 590080 560898
rect 589460 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 590080 525454
rect 589460 525134 590080 525218
rect 589460 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 590080 525134
rect 589460 489454 590080 524898
rect 589460 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 590080 489454
rect 589460 489134 590080 489218
rect 589460 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 590080 489134
rect 589460 453454 590080 488898
rect 589460 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 590080 453454
rect 589460 453134 590080 453218
rect 589460 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 590080 453134
rect 589460 417454 590080 452898
rect 589460 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 590080 417454
rect 589460 417134 590080 417218
rect 589460 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 590080 417134
rect 589460 381454 590080 416898
rect 589460 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 590080 381454
rect 589460 381134 590080 381218
rect 589460 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 590080 381134
rect 589460 345454 590080 380898
rect 589460 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 590080 345454
rect 589460 345134 590080 345218
rect 589460 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 590080 345134
rect 589460 309454 590080 344898
rect 589460 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 590080 309454
rect 589460 309134 590080 309218
rect 589460 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 590080 309134
rect 589460 273454 590080 308898
rect 589460 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 590080 273454
rect 589460 273134 590080 273218
rect 589460 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 590080 273134
rect 589460 237454 590080 272898
rect 589460 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 590080 237454
rect 589460 237134 590080 237218
rect 589460 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 590080 237134
rect 589460 201454 590080 236898
rect 589460 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 590080 201454
rect 589460 201134 590080 201218
rect 589460 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 590080 201134
rect 589460 165454 590080 200898
rect 589460 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 590080 165454
rect 589460 165134 590080 165218
rect 589460 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 590080 165134
rect 589460 129454 590080 164898
rect 589460 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 590080 129454
rect 589460 129134 590080 129218
rect 589460 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 590080 129134
rect 589460 93454 590080 128898
rect 589460 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 590080 93454
rect 589460 93134 590080 93218
rect 589460 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 590080 93134
rect 589460 57454 590080 92898
rect 589460 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 590080 57454
rect 589460 57134 590080 57218
rect 589460 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 590080 57134
rect 589460 21454 590080 56898
rect 589460 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 590080 21454
rect 589460 21134 590080 21218
rect 589460 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 590080 21134
rect 589460 -4496 590080 20898
rect 589460 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect 589460 -4816 590080 -4732
rect 589460 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect 589460 -5084 590080 -5052
rect 590420 673954 591040 709392
rect 590420 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 591040 673954
rect 590420 673634 591040 673718
rect 590420 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 591040 673634
rect 590420 637954 591040 673398
rect 590420 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 591040 637954
rect 590420 637634 591040 637718
rect 590420 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 591040 637634
rect 590420 601954 591040 637398
rect 590420 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 591040 601954
rect 590420 601634 591040 601718
rect 590420 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 591040 601634
rect 590420 565954 591040 601398
rect 590420 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 591040 565954
rect 590420 565634 591040 565718
rect 590420 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 591040 565634
rect 590420 529954 591040 565398
rect 590420 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 591040 529954
rect 590420 529634 591040 529718
rect 590420 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 591040 529634
rect 590420 493954 591040 529398
rect 590420 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 591040 493954
rect 590420 493634 591040 493718
rect 590420 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 591040 493634
rect 590420 457954 591040 493398
rect 590420 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 591040 457954
rect 590420 457634 591040 457718
rect 590420 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 591040 457634
rect 590420 421954 591040 457398
rect 590420 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 591040 421954
rect 590420 421634 591040 421718
rect 590420 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 591040 421634
rect 590420 385954 591040 421398
rect 590420 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 591040 385954
rect 590420 385634 591040 385718
rect 590420 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 591040 385634
rect 590420 349954 591040 385398
rect 590420 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 591040 349954
rect 590420 349634 591040 349718
rect 590420 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 591040 349634
rect 590420 313954 591040 349398
rect 590420 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 591040 313954
rect 590420 313634 591040 313718
rect 590420 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 591040 313634
rect 590420 277954 591040 313398
rect 590420 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 591040 277954
rect 590420 277634 591040 277718
rect 590420 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 591040 277634
rect 590420 241954 591040 277398
rect 590420 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 591040 241954
rect 590420 241634 591040 241718
rect 590420 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 591040 241634
rect 590420 205954 591040 241398
rect 590420 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 591040 205954
rect 590420 205634 591040 205718
rect 590420 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 591040 205634
rect 590420 169954 591040 205398
rect 590420 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 591040 169954
rect 590420 169634 591040 169718
rect 590420 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 591040 169634
rect 590420 133954 591040 169398
rect 590420 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 591040 133954
rect 590420 133634 591040 133718
rect 590420 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 591040 133634
rect 590420 97954 591040 133398
rect 590420 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 591040 97954
rect 590420 97634 591040 97718
rect 590420 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 591040 97634
rect 590420 61954 591040 97398
rect 590420 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 591040 61954
rect 590420 61634 591040 61718
rect 590420 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 591040 61634
rect 590420 25954 591040 61398
rect 590420 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 591040 25954
rect 590420 25634 591040 25718
rect 590420 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 591040 25634
rect 590420 -5456 591040 25398
rect 590420 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect 590420 -5776 591040 -5692
rect 590420 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect 590420 -6044 591040 -6012
rect 591380 678454 592000 710352
rect 591380 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592000 678454
rect 591380 678134 592000 678218
rect 591380 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592000 678134
rect 591380 642454 592000 677898
rect 591380 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592000 642454
rect 591380 642134 592000 642218
rect 591380 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592000 642134
rect 591380 606454 592000 641898
rect 591380 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592000 606454
rect 591380 606134 592000 606218
rect 591380 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592000 606134
rect 591380 570454 592000 605898
rect 591380 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592000 570454
rect 591380 570134 592000 570218
rect 591380 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592000 570134
rect 591380 534454 592000 569898
rect 591380 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592000 534454
rect 591380 534134 592000 534218
rect 591380 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592000 534134
rect 591380 498454 592000 533898
rect 591380 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592000 498454
rect 591380 498134 592000 498218
rect 591380 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592000 498134
rect 591380 462454 592000 497898
rect 591380 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592000 462454
rect 591380 462134 592000 462218
rect 591380 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592000 462134
rect 591380 426454 592000 461898
rect 591380 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592000 426454
rect 591380 426134 592000 426218
rect 591380 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592000 426134
rect 591380 390454 592000 425898
rect 591380 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592000 390454
rect 591380 390134 592000 390218
rect 591380 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592000 390134
rect 591380 354454 592000 389898
rect 591380 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592000 354454
rect 591380 354134 592000 354218
rect 591380 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592000 354134
rect 591380 318454 592000 353898
rect 591380 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592000 318454
rect 591380 318134 592000 318218
rect 591380 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592000 318134
rect 591380 282454 592000 317898
rect 591380 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592000 282454
rect 591380 282134 592000 282218
rect 591380 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592000 282134
rect 591380 246454 592000 281898
rect 591380 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592000 246454
rect 591380 246134 592000 246218
rect 591380 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592000 246134
rect 591380 210454 592000 245898
rect 591380 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592000 210454
rect 591380 210134 592000 210218
rect 591380 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592000 210134
rect 591380 174454 592000 209898
rect 591380 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592000 174454
rect 591380 174134 592000 174218
rect 591380 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592000 174134
rect 591380 138454 592000 173898
rect 591380 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592000 138454
rect 591380 138134 592000 138218
rect 591380 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592000 138134
rect 591380 102454 592000 137898
rect 591380 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592000 102454
rect 591380 102134 592000 102218
rect 591380 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592000 102134
rect 591380 66454 592000 101898
rect 591380 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592000 66454
rect 591380 66134 592000 66218
rect 591380 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592000 66134
rect 591380 30454 592000 65898
rect 591380 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592000 30454
rect 591380 30134 592000 30218
rect 591380 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592000 30134
rect 591380 -6416 592000 29898
rect 591380 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect 591380 -6736 592000 -6652
rect 591380 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect 591380 -7004 592000 -6972
rect 592340 682954 592960 711312
rect 592340 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect 592340 682634 592960 682718
rect 592340 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect 592340 646954 592960 682398
rect 592340 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect 592340 646634 592960 646718
rect 592340 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect 592340 610954 592960 646398
rect 592340 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect 592340 610634 592960 610718
rect 592340 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect 592340 574954 592960 610398
rect 592340 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect 592340 574634 592960 574718
rect 592340 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect 592340 538954 592960 574398
rect 592340 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect 592340 538634 592960 538718
rect 592340 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect 592340 502954 592960 538398
rect 592340 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect 592340 502634 592960 502718
rect 592340 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect 592340 466954 592960 502398
rect 592340 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect 592340 466634 592960 466718
rect 592340 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect 592340 430954 592960 466398
rect 592340 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect 592340 430634 592960 430718
rect 592340 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect 592340 394954 592960 430398
rect 592340 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect 592340 394634 592960 394718
rect 592340 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect 592340 358954 592960 394398
rect 592340 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect 592340 358634 592960 358718
rect 592340 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect 592340 322954 592960 358398
rect 592340 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect 592340 322634 592960 322718
rect 592340 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect 592340 286954 592960 322398
rect 592340 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect 592340 286634 592960 286718
rect 592340 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect 592340 250954 592960 286398
rect 592340 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect 592340 250634 592960 250718
rect 592340 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect 592340 214954 592960 250398
rect 592340 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect 592340 214634 592960 214718
rect 592340 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect 592340 178954 592960 214398
rect 592340 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect 592340 178634 592960 178718
rect 592340 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect 592340 142954 592960 178398
rect 592340 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect 592340 142634 592960 142718
rect 592340 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect 592340 106954 592960 142398
rect 592340 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect 592340 106634 592960 106718
rect 592340 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect 592340 70954 592960 106398
rect 592340 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect 592340 70634 592960 70718
rect 592340 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect 592340 34954 592960 70398
rect 592340 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect 592340 34634 592960 34718
rect 592340 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect 592340 -7376 592960 34398
rect 592340 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect 592340 -7696 592960 -7612
rect 592340 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect 592340 -7964 592960 -7932
<< via4 >>
rect -9004 711632 -8768 711868
rect -8684 711632 -8448 711868
rect -9004 711312 -8768 711548
rect -8684 711312 -8448 711548
rect -9004 682718 -8768 682954
rect -8684 682718 -8448 682954
rect -9004 682398 -8768 682634
rect -8684 682398 -8448 682634
rect -9004 646718 -8768 646954
rect -8684 646718 -8448 646954
rect -9004 646398 -8768 646634
rect -8684 646398 -8448 646634
rect -9004 610718 -8768 610954
rect -8684 610718 -8448 610954
rect -9004 610398 -8768 610634
rect -8684 610398 -8448 610634
rect -9004 574718 -8768 574954
rect -8684 574718 -8448 574954
rect -9004 574398 -8768 574634
rect -8684 574398 -8448 574634
rect -9004 538718 -8768 538954
rect -8684 538718 -8448 538954
rect -9004 538398 -8768 538634
rect -8684 538398 -8448 538634
rect -9004 502718 -8768 502954
rect -8684 502718 -8448 502954
rect -9004 502398 -8768 502634
rect -8684 502398 -8448 502634
rect -9004 466718 -8768 466954
rect -8684 466718 -8448 466954
rect -9004 466398 -8768 466634
rect -8684 466398 -8448 466634
rect -9004 430718 -8768 430954
rect -8684 430718 -8448 430954
rect -9004 430398 -8768 430634
rect -8684 430398 -8448 430634
rect -9004 394718 -8768 394954
rect -8684 394718 -8448 394954
rect -9004 394398 -8768 394634
rect -8684 394398 -8448 394634
rect -9004 358718 -8768 358954
rect -8684 358718 -8448 358954
rect -9004 358398 -8768 358634
rect -8684 358398 -8448 358634
rect -9004 322718 -8768 322954
rect -8684 322718 -8448 322954
rect -9004 322398 -8768 322634
rect -8684 322398 -8448 322634
rect -9004 286718 -8768 286954
rect -8684 286718 -8448 286954
rect -9004 286398 -8768 286634
rect -8684 286398 -8448 286634
rect -9004 250718 -8768 250954
rect -8684 250718 -8448 250954
rect -9004 250398 -8768 250634
rect -8684 250398 -8448 250634
rect -9004 214718 -8768 214954
rect -8684 214718 -8448 214954
rect -9004 214398 -8768 214634
rect -8684 214398 -8448 214634
rect -9004 178718 -8768 178954
rect -8684 178718 -8448 178954
rect -9004 178398 -8768 178634
rect -8684 178398 -8448 178634
rect -9004 142718 -8768 142954
rect -8684 142718 -8448 142954
rect -9004 142398 -8768 142634
rect -8684 142398 -8448 142634
rect -9004 106718 -8768 106954
rect -8684 106718 -8448 106954
rect -9004 106398 -8768 106634
rect -8684 106398 -8448 106634
rect -9004 70718 -8768 70954
rect -8684 70718 -8448 70954
rect -9004 70398 -8768 70634
rect -8684 70398 -8448 70634
rect -9004 34718 -8768 34954
rect -8684 34718 -8448 34954
rect -9004 34398 -8768 34634
rect -8684 34398 -8448 34634
rect -8044 710672 -7808 710908
rect -7724 710672 -7488 710908
rect -8044 710352 -7808 710588
rect -7724 710352 -7488 710588
rect -8044 678218 -7808 678454
rect -7724 678218 -7488 678454
rect -8044 677898 -7808 678134
rect -7724 677898 -7488 678134
rect -8044 642218 -7808 642454
rect -7724 642218 -7488 642454
rect -8044 641898 -7808 642134
rect -7724 641898 -7488 642134
rect -8044 606218 -7808 606454
rect -7724 606218 -7488 606454
rect -8044 605898 -7808 606134
rect -7724 605898 -7488 606134
rect -8044 570218 -7808 570454
rect -7724 570218 -7488 570454
rect -8044 569898 -7808 570134
rect -7724 569898 -7488 570134
rect -8044 534218 -7808 534454
rect -7724 534218 -7488 534454
rect -8044 533898 -7808 534134
rect -7724 533898 -7488 534134
rect -8044 498218 -7808 498454
rect -7724 498218 -7488 498454
rect -8044 497898 -7808 498134
rect -7724 497898 -7488 498134
rect -8044 462218 -7808 462454
rect -7724 462218 -7488 462454
rect -8044 461898 -7808 462134
rect -7724 461898 -7488 462134
rect -8044 426218 -7808 426454
rect -7724 426218 -7488 426454
rect -8044 425898 -7808 426134
rect -7724 425898 -7488 426134
rect -8044 390218 -7808 390454
rect -7724 390218 -7488 390454
rect -8044 389898 -7808 390134
rect -7724 389898 -7488 390134
rect -8044 354218 -7808 354454
rect -7724 354218 -7488 354454
rect -8044 353898 -7808 354134
rect -7724 353898 -7488 354134
rect -8044 318218 -7808 318454
rect -7724 318218 -7488 318454
rect -8044 317898 -7808 318134
rect -7724 317898 -7488 318134
rect -8044 282218 -7808 282454
rect -7724 282218 -7488 282454
rect -8044 281898 -7808 282134
rect -7724 281898 -7488 282134
rect -8044 246218 -7808 246454
rect -7724 246218 -7488 246454
rect -8044 245898 -7808 246134
rect -7724 245898 -7488 246134
rect -8044 210218 -7808 210454
rect -7724 210218 -7488 210454
rect -8044 209898 -7808 210134
rect -7724 209898 -7488 210134
rect -8044 174218 -7808 174454
rect -7724 174218 -7488 174454
rect -8044 173898 -7808 174134
rect -7724 173898 -7488 174134
rect -8044 138218 -7808 138454
rect -7724 138218 -7488 138454
rect -8044 137898 -7808 138134
rect -7724 137898 -7488 138134
rect -8044 102218 -7808 102454
rect -7724 102218 -7488 102454
rect -8044 101898 -7808 102134
rect -7724 101898 -7488 102134
rect -8044 66218 -7808 66454
rect -7724 66218 -7488 66454
rect -8044 65898 -7808 66134
rect -7724 65898 -7488 66134
rect -8044 30218 -7808 30454
rect -7724 30218 -7488 30454
rect -8044 29898 -7808 30134
rect -7724 29898 -7488 30134
rect -7084 709712 -6848 709948
rect -6764 709712 -6528 709948
rect -7084 709392 -6848 709628
rect -6764 709392 -6528 709628
rect -7084 673718 -6848 673954
rect -6764 673718 -6528 673954
rect -7084 673398 -6848 673634
rect -6764 673398 -6528 673634
rect -7084 637718 -6848 637954
rect -6764 637718 -6528 637954
rect -7084 637398 -6848 637634
rect -6764 637398 -6528 637634
rect -7084 601718 -6848 601954
rect -6764 601718 -6528 601954
rect -7084 601398 -6848 601634
rect -6764 601398 -6528 601634
rect -7084 565718 -6848 565954
rect -6764 565718 -6528 565954
rect -7084 565398 -6848 565634
rect -6764 565398 -6528 565634
rect -7084 529718 -6848 529954
rect -6764 529718 -6528 529954
rect -7084 529398 -6848 529634
rect -6764 529398 -6528 529634
rect -7084 493718 -6848 493954
rect -6764 493718 -6528 493954
rect -7084 493398 -6848 493634
rect -6764 493398 -6528 493634
rect -7084 457718 -6848 457954
rect -6764 457718 -6528 457954
rect -7084 457398 -6848 457634
rect -6764 457398 -6528 457634
rect -7084 421718 -6848 421954
rect -6764 421718 -6528 421954
rect -7084 421398 -6848 421634
rect -6764 421398 -6528 421634
rect -7084 385718 -6848 385954
rect -6764 385718 -6528 385954
rect -7084 385398 -6848 385634
rect -6764 385398 -6528 385634
rect -7084 349718 -6848 349954
rect -6764 349718 -6528 349954
rect -7084 349398 -6848 349634
rect -6764 349398 -6528 349634
rect -7084 313718 -6848 313954
rect -6764 313718 -6528 313954
rect -7084 313398 -6848 313634
rect -6764 313398 -6528 313634
rect -7084 277718 -6848 277954
rect -6764 277718 -6528 277954
rect -7084 277398 -6848 277634
rect -6764 277398 -6528 277634
rect -7084 241718 -6848 241954
rect -6764 241718 -6528 241954
rect -7084 241398 -6848 241634
rect -6764 241398 -6528 241634
rect -7084 205718 -6848 205954
rect -6764 205718 -6528 205954
rect -7084 205398 -6848 205634
rect -6764 205398 -6528 205634
rect -7084 169718 -6848 169954
rect -6764 169718 -6528 169954
rect -7084 169398 -6848 169634
rect -6764 169398 -6528 169634
rect -7084 133718 -6848 133954
rect -6764 133718 -6528 133954
rect -7084 133398 -6848 133634
rect -6764 133398 -6528 133634
rect -7084 97718 -6848 97954
rect -6764 97718 -6528 97954
rect -7084 97398 -6848 97634
rect -6764 97398 -6528 97634
rect -7084 61718 -6848 61954
rect -6764 61718 -6528 61954
rect -7084 61398 -6848 61634
rect -6764 61398 -6528 61634
rect -7084 25718 -6848 25954
rect -6764 25718 -6528 25954
rect -7084 25398 -6848 25634
rect -6764 25398 -6528 25634
rect -6124 708752 -5888 708988
rect -5804 708752 -5568 708988
rect -6124 708432 -5888 708668
rect -5804 708432 -5568 708668
rect -6124 669218 -5888 669454
rect -5804 669218 -5568 669454
rect -6124 668898 -5888 669134
rect -5804 668898 -5568 669134
rect -6124 633218 -5888 633454
rect -5804 633218 -5568 633454
rect -6124 632898 -5888 633134
rect -5804 632898 -5568 633134
rect -6124 597218 -5888 597454
rect -5804 597218 -5568 597454
rect -6124 596898 -5888 597134
rect -5804 596898 -5568 597134
rect -6124 561218 -5888 561454
rect -5804 561218 -5568 561454
rect -6124 560898 -5888 561134
rect -5804 560898 -5568 561134
rect -6124 525218 -5888 525454
rect -5804 525218 -5568 525454
rect -6124 524898 -5888 525134
rect -5804 524898 -5568 525134
rect -6124 489218 -5888 489454
rect -5804 489218 -5568 489454
rect -6124 488898 -5888 489134
rect -5804 488898 -5568 489134
rect -6124 453218 -5888 453454
rect -5804 453218 -5568 453454
rect -6124 452898 -5888 453134
rect -5804 452898 -5568 453134
rect -6124 417218 -5888 417454
rect -5804 417218 -5568 417454
rect -6124 416898 -5888 417134
rect -5804 416898 -5568 417134
rect -6124 381218 -5888 381454
rect -5804 381218 -5568 381454
rect -6124 380898 -5888 381134
rect -5804 380898 -5568 381134
rect -6124 345218 -5888 345454
rect -5804 345218 -5568 345454
rect -6124 344898 -5888 345134
rect -5804 344898 -5568 345134
rect -6124 309218 -5888 309454
rect -5804 309218 -5568 309454
rect -6124 308898 -5888 309134
rect -5804 308898 -5568 309134
rect -6124 273218 -5888 273454
rect -5804 273218 -5568 273454
rect -6124 272898 -5888 273134
rect -5804 272898 -5568 273134
rect -6124 237218 -5888 237454
rect -5804 237218 -5568 237454
rect -6124 236898 -5888 237134
rect -5804 236898 -5568 237134
rect -6124 201218 -5888 201454
rect -5804 201218 -5568 201454
rect -6124 200898 -5888 201134
rect -5804 200898 -5568 201134
rect -6124 165218 -5888 165454
rect -5804 165218 -5568 165454
rect -6124 164898 -5888 165134
rect -5804 164898 -5568 165134
rect -6124 129218 -5888 129454
rect -5804 129218 -5568 129454
rect -6124 128898 -5888 129134
rect -5804 128898 -5568 129134
rect -6124 93218 -5888 93454
rect -5804 93218 -5568 93454
rect -6124 92898 -5888 93134
rect -5804 92898 -5568 93134
rect -6124 57218 -5888 57454
rect -5804 57218 -5568 57454
rect -6124 56898 -5888 57134
rect -5804 56898 -5568 57134
rect -6124 21218 -5888 21454
rect -5804 21218 -5568 21454
rect -6124 20898 -5888 21134
rect -5804 20898 -5568 21134
rect -5164 707792 -4928 708028
rect -4844 707792 -4608 708028
rect -5164 707472 -4928 707708
rect -4844 707472 -4608 707708
rect -5164 700718 -4928 700954
rect -4844 700718 -4608 700954
rect -5164 700398 -4928 700634
rect -4844 700398 -4608 700634
rect -5164 664718 -4928 664954
rect -4844 664718 -4608 664954
rect -5164 664398 -4928 664634
rect -4844 664398 -4608 664634
rect -5164 628718 -4928 628954
rect -4844 628718 -4608 628954
rect -5164 628398 -4928 628634
rect -4844 628398 -4608 628634
rect -5164 592718 -4928 592954
rect -4844 592718 -4608 592954
rect -5164 592398 -4928 592634
rect -4844 592398 -4608 592634
rect -5164 556718 -4928 556954
rect -4844 556718 -4608 556954
rect -5164 556398 -4928 556634
rect -4844 556398 -4608 556634
rect -5164 520718 -4928 520954
rect -4844 520718 -4608 520954
rect -5164 520398 -4928 520634
rect -4844 520398 -4608 520634
rect -5164 484718 -4928 484954
rect -4844 484718 -4608 484954
rect -5164 484398 -4928 484634
rect -4844 484398 -4608 484634
rect -5164 448718 -4928 448954
rect -4844 448718 -4608 448954
rect -5164 448398 -4928 448634
rect -4844 448398 -4608 448634
rect -5164 412718 -4928 412954
rect -4844 412718 -4608 412954
rect -5164 412398 -4928 412634
rect -4844 412398 -4608 412634
rect -5164 376718 -4928 376954
rect -4844 376718 -4608 376954
rect -5164 376398 -4928 376634
rect -4844 376398 -4608 376634
rect -5164 340718 -4928 340954
rect -4844 340718 -4608 340954
rect -5164 340398 -4928 340634
rect -4844 340398 -4608 340634
rect -5164 304718 -4928 304954
rect -4844 304718 -4608 304954
rect -5164 304398 -4928 304634
rect -4844 304398 -4608 304634
rect -5164 268718 -4928 268954
rect -4844 268718 -4608 268954
rect -5164 268398 -4928 268634
rect -4844 268398 -4608 268634
rect -5164 232718 -4928 232954
rect -4844 232718 -4608 232954
rect -5164 232398 -4928 232634
rect -4844 232398 -4608 232634
rect -5164 196718 -4928 196954
rect -4844 196718 -4608 196954
rect -5164 196398 -4928 196634
rect -4844 196398 -4608 196634
rect -5164 160718 -4928 160954
rect -4844 160718 -4608 160954
rect -5164 160398 -4928 160634
rect -4844 160398 -4608 160634
rect -5164 124718 -4928 124954
rect -4844 124718 -4608 124954
rect -5164 124398 -4928 124634
rect -4844 124398 -4608 124634
rect -5164 88718 -4928 88954
rect -4844 88718 -4608 88954
rect -5164 88398 -4928 88634
rect -4844 88398 -4608 88634
rect -5164 52718 -4928 52954
rect -4844 52718 -4608 52954
rect -5164 52398 -4928 52634
rect -4844 52398 -4608 52634
rect -5164 16718 -4928 16954
rect -4844 16718 -4608 16954
rect -5164 16398 -4928 16634
rect -4844 16398 -4608 16634
rect -4204 706832 -3968 707068
rect -3884 706832 -3648 707068
rect -4204 706512 -3968 706748
rect -3884 706512 -3648 706748
rect -4204 696218 -3968 696454
rect -3884 696218 -3648 696454
rect -4204 695898 -3968 696134
rect -3884 695898 -3648 696134
rect -4204 660218 -3968 660454
rect -3884 660218 -3648 660454
rect -4204 659898 -3968 660134
rect -3884 659898 -3648 660134
rect -4204 624218 -3968 624454
rect -3884 624218 -3648 624454
rect -4204 623898 -3968 624134
rect -3884 623898 -3648 624134
rect -4204 588218 -3968 588454
rect -3884 588218 -3648 588454
rect -4204 587898 -3968 588134
rect -3884 587898 -3648 588134
rect -4204 552218 -3968 552454
rect -3884 552218 -3648 552454
rect -4204 551898 -3968 552134
rect -3884 551898 -3648 552134
rect -4204 516218 -3968 516454
rect -3884 516218 -3648 516454
rect -4204 515898 -3968 516134
rect -3884 515898 -3648 516134
rect -4204 480218 -3968 480454
rect -3884 480218 -3648 480454
rect -4204 479898 -3968 480134
rect -3884 479898 -3648 480134
rect -4204 444218 -3968 444454
rect -3884 444218 -3648 444454
rect -4204 443898 -3968 444134
rect -3884 443898 -3648 444134
rect -4204 408218 -3968 408454
rect -3884 408218 -3648 408454
rect -4204 407898 -3968 408134
rect -3884 407898 -3648 408134
rect -4204 372218 -3968 372454
rect -3884 372218 -3648 372454
rect -4204 371898 -3968 372134
rect -3884 371898 -3648 372134
rect -4204 336218 -3968 336454
rect -3884 336218 -3648 336454
rect -4204 335898 -3968 336134
rect -3884 335898 -3648 336134
rect -4204 300218 -3968 300454
rect -3884 300218 -3648 300454
rect -4204 299898 -3968 300134
rect -3884 299898 -3648 300134
rect -4204 264218 -3968 264454
rect -3884 264218 -3648 264454
rect -4204 263898 -3968 264134
rect -3884 263898 -3648 264134
rect -4204 228218 -3968 228454
rect -3884 228218 -3648 228454
rect -4204 227898 -3968 228134
rect -3884 227898 -3648 228134
rect -4204 192218 -3968 192454
rect -3884 192218 -3648 192454
rect -4204 191898 -3968 192134
rect -3884 191898 -3648 192134
rect -4204 156218 -3968 156454
rect -3884 156218 -3648 156454
rect -4204 155898 -3968 156134
rect -3884 155898 -3648 156134
rect -4204 120218 -3968 120454
rect -3884 120218 -3648 120454
rect -4204 119898 -3968 120134
rect -3884 119898 -3648 120134
rect -4204 84218 -3968 84454
rect -3884 84218 -3648 84454
rect -4204 83898 -3968 84134
rect -3884 83898 -3648 84134
rect -4204 48218 -3968 48454
rect -3884 48218 -3648 48454
rect -4204 47898 -3968 48134
rect -3884 47898 -3648 48134
rect -4204 12218 -3968 12454
rect -3884 12218 -3648 12454
rect -4204 11898 -3968 12134
rect -3884 11898 -3648 12134
rect -3244 705872 -3008 706108
rect -2924 705872 -2688 706108
rect -3244 705552 -3008 705788
rect -2924 705552 -2688 705788
rect -3244 691718 -3008 691954
rect -2924 691718 -2688 691954
rect -3244 691398 -3008 691634
rect -2924 691398 -2688 691634
rect -3244 655718 -3008 655954
rect -2924 655718 -2688 655954
rect -3244 655398 -3008 655634
rect -2924 655398 -2688 655634
rect -3244 619718 -3008 619954
rect -2924 619718 -2688 619954
rect -3244 619398 -3008 619634
rect -2924 619398 -2688 619634
rect -3244 583718 -3008 583954
rect -2924 583718 -2688 583954
rect -3244 583398 -3008 583634
rect -2924 583398 -2688 583634
rect -3244 547718 -3008 547954
rect -2924 547718 -2688 547954
rect -3244 547398 -3008 547634
rect -2924 547398 -2688 547634
rect -3244 511718 -3008 511954
rect -2924 511718 -2688 511954
rect -3244 511398 -3008 511634
rect -2924 511398 -2688 511634
rect -3244 475718 -3008 475954
rect -2924 475718 -2688 475954
rect -3244 475398 -3008 475634
rect -2924 475398 -2688 475634
rect -3244 439718 -3008 439954
rect -2924 439718 -2688 439954
rect -3244 439398 -3008 439634
rect -2924 439398 -2688 439634
rect -3244 403718 -3008 403954
rect -2924 403718 -2688 403954
rect -3244 403398 -3008 403634
rect -2924 403398 -2688 403634
rect -3244 367718 -3008 367954
rect -2924 367718 -2688 367954
rect -3244 367398 -3008 367634
rect -2924 367398 -2688 367634
rect -3244 331718 -3008 331954
rect -2924 331718 -2688 331954
rect -3244 331398 -3008 331634
rect -2924 331398 -2688 331634
rect -3244 295718 -3008 295954
rect -2924 295718 -2688 295954
rect -3244 295398 -3008 295634
rect -2924 295398 -2688 295634
rect -3244 259718 -3008 259954
rect -2924 259718 -2688 259954
rect -3244 259398 -3008 259634
rect -2924 259398 -2688 259634
rect -3244 223718 -3008 223954
rect -2924 223718 -2688 223954
rect -3244 223398 -3008 223634
rect -2924 223398 -2688 223634
rect -3244 187718 -3008 187954
rect -2924 187718 -2688 187954
rect -3244 187398 -3008 187634
rect -2924 187398 -2688 187634
rect -3244 151718 -3008 151954
rect -2924 151718 -2688 151954
rect -3244 151398 -3008 151634
rect -2924 151398 -2688 151634
rect -3244 115718 -3008 115954
rect -2924 115718 -2688 115954
rect -3244 115398 -3008 115634
rect -2924 115398 -2688 115634
rect -3244 79718 -3008 79954
rect -2924 79718 -2688 79954
rect -3244 79398 -3008 79634
rect -2924 79398 -2688 79634
rect -3244 43718 -3008 43954
rect -2924 43718 -2688 43954
rect -3244 43398 -3008 43634
rect -2924 43398 -2688 43634
rect -3244 7718 -3008 7954
rect -2924 7718 -2688 7954
rect -3244 7398 -3008 7634
rect -2924 7398 -2688 7634
rect -2284 704912 -2048 705148
rect -1964 704912 -1728 705148
rect -2284 704592 -2048 704828
rect -1964 704592 -1728 704828
rect -2284 687218 -2048 687454
rect -1964 687218 -1728 687454
rect -2284 686898 -2048 687134
rect -1964 686898 -1728 687134
rect -2284 651218 -2048 651454
rect -1964 651218 -1728 651454
rect -2284 650898 -2048 651134
rect -1964 650898 -1728 651134
rect -2284 615218 -2048 615454
rect -1964 615218 -1728 615454
rect -2284 614898 -2048 615134
rect -1964 614898 -1728 615134
rect -2284 579218 -2048 579454
rect -1964 579218 -1728 579454
rect -2284 578898 -2048 579134
rect -1964 578898 -1728 579134
rect -2284 543218 -2048 543454
rect -1964 543218 -1728 543454
rect -2284 542898 -2048 543134
rect -1964 542898 -1728 543134
rect -2284 507218 -2048 507454
rect -1964 507218 -1728 507454
rect -2284 506898 -2048 507134
rect -1964 506898 -1728 507134
rect -2284 471218 -2048 471454
rect -1964 471218 -1728 471454
rect -2284 470898 -2048 471134
rect -1964 470898 -1728 471134
rect -2284 435218 -2048 435454
rect -1964 435218 -1728 435454
rect -2284 434898 -2048 435134
rect -1964 434898 -1728 435134
rect -2284 399218 -2048 399454
rect -1964 399218 -1728 399454
rect -2284 398898 -2048 399134
rect -1964 398898 -1728 399134
rect -2284 363218 -2048 363454
rect -1964 363218 -1728 363454
rect -2284 362898 -2048 363134
rect -1964 362898 -1728 363134
rect -2284 327218 -2048 327454
rect -1964 327218 -1728 327454
rect -2284 326898 -2048 327134
rect -1964 326898 -1728 327134
rect -2284 291218 -2048 291454
rect -1964 291218 -1728 291454
rect -2284 290898 -2048 291134
rect -1964 290898 -1728 291134
rect -2284 255218 -2048 255454
rect -1964 255218 -1728 255454
rect -2284 254898 -2048 255134
rect -1964 254898 -1728 255134
rect -2284 219218 -2048 219454
rect -1964 219218 -1728 219454
rect -2284 218898 -2048 219134
rect -1964 218898 -1728 219134
rect -2284 183218 -2048 183454
rect -1964 183218 -1728 183454
rect -2284 182898 -2048 183134
rect -1964 182898 -1728 183134
rect -2284 147218 -2048 147454
rect -1964 147218 -1728 147454
rect -2284 146898 -2048 147134
rect -1964 146898 -1728 147134
rect -2284 111218 -2048 111454
rect -1964 111218 -1728 111454
rect -2284 110898 -2048 111134
rect -1964 110898 -1728 111134
rect -2284 75218 -2048 75454
rect -1964 75218 -1728 75454
rect -2284 74898 -2048 75134
rect -1964 74898 -1728 75134
rect -2284 39218 -2048 39454
rect -1964 39218 -1728 39454
rect -2284 38898 -2048 39134
rect -1964 38898 -1728 39134
rect -2284 3218 -2048 3454
rect -1964 3218 -1728 3454
rect -2284 2898 -2048 3134
rect -1964 2898 -1728 3134
rect -2284 -892 -2048 -656
rect -1964 -892 -1728 -656
rect -2284 -1212 -2048 -976
rect -1964 -1212 -1728 -976
rect 1826 704912 2062 705148
rect 2146 704912 2382 705148
rect 1826 704592 2062 704828
rect 2146 704592 2382 704828
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -892 2062 -656
rect 2146 -892 2382 -656
rect 1826 -1212 2062 -976
rect 2146 -1212 2382 -976
rect -3244 -1852 -3008 -1616
rect -2924 -1852 -2688 -1616
rect -3244 -2172 -3008 -1936
rect -2924 -2172 -2688 -1936
rect -4204 -2812 -3968 -2576
rect -3884 -2812 -3648 -2576
rect -4204 -3132 -3968 -2896
rect -3884 -3132 -3648 -2896
rect -5164 -3772 -4928 -3536
rect -4844 -3772 -4608 -3536
rect -5164 -4092 -4928 -3856
rect -4844 -4092 -4608 -3856
rect -6124 -4732 -5888 -4496
rect -5804 -4732 -5568 -4496
rect -6124 -5052 -5888 -4816
rect -5804 -5052 -5568 -4816
rect -7084 -5692 -6848 -5456
rect -6764 -5692 -6528 -5456
rect -7084 -6012 -6848 -5776
rect -6764 -6012 -6528 -5776
rect -8044 -6652 -7808 -6416
rect -7724 -6652 -7488 -6416
rect -8044 -6972 -7808 -6736
rect -7724 -6972 -7488 -6736
rect -9004 -7612 -8768 -7376
rect -8684 -7612 -8448 -7376
rect -9004 -7932 -8768 -7696
rect -8684 -7932 -8448 -7696
rect 6326 705872 6562 706108
rect 6646 705872 6882 706108
rect 6326 705552 6562 705788
rect 6646 705552 6882 705788
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1852 6562 -1616
rect 6646 -1852 6882 -1616
rect 6326 -2172 6562 -1936
rect 6646 -2172 6882 -1936
rect 10826 706832 11062 707068
rect 11146 706832 11382 707068
rect 10826 706512 11062 706748
rect 11146 706512 11382 706748
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2812 11062 -2576
rect 11146 -2812 11382 -2576
rect 10826 -3132 11062 -2896
rect 11146 -3132 11382 -2896
rect 15326 707792 15562 708028
rect 15646 707792 15882 708028
rect 15326 707472 15562 707708
rect 15646 707472 15882 707708
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3772 15562 -3536
rect 15646 -3772 15882 -3536
rect 15326 -4092 15562 -3856
rect 15646 -4092 15882 -3856
rect 19826 708752 20062 708988
rect 20146 708752 20382 708988
rect 19826 708432 20062 708668
rect 20146 708432 20382 708668
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4732 20062 -4496
rect 20146 -4732 20382 -4496
rect 19826 -5052 20062 -4816
rect 20146 -5052 20382 -4816
rect 24326 709712 24562 709948
rect 24646 709712 24882 709948
rect 24326 709392 24562 709628
rect 24646 709392 24882 709628
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5692 24562 -5456
rect 24646 -5692 24882 -5456
rect 24326 -6012 24562 -5776
rect 24646 -6012 24882 -5776
rect 28826 710672 29062 710908
rect 29146 710672 29382 710908
rect 28826 710352 29062 710588
rect 29146 710352 29382 710588
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6652 29062 -6416
rect 29146 -6652 29382 -6416
rect 28826 -6972 29062 -6736
rect 29146 -6972 29382 -6736
rect 33326 711632 33562 711868
rect 33646 711632 33882 711868
rect 33326 711312 33562 711548
rect 33646 711312 33882 711548
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7612 33562 -7376
rect 33646 -7612 33882 -7376
rect 33326 -7932 33562 -7696
rect 33646 -7932 33882 -7696
rect 37826 704912 38062 705148
rect 38146 704912 38382 705148
rect 37826 704592 38062 704828
rect 38146 704592 38382 704828
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -892 38062 -656
rect 38146 -892 38382 -656
rect 37826 -1212 38062 -976
rect 38146 -1212 38382 -976
rect 42326 705872 42562 706108
rect 42646 705872 42882 706108
rect 42326 705552 42562 705788
rect 42646 705552 42882 705788
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1852 42562 -1616
rect 42646 -1852 42882 -1616
rect 42326 -2172 42562 -1936
rect 42646 -2172 42882 -1936
rect 46826 706832 47062 707068
rect 47146 706832 47382 707068
rect 46826 706512 47062 706748
rect 47146 706512 47382 706748
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2812 47062 -2576
rect 47146 -2812 47382 -2576
rect 46826 -3132 47062 -2896
rect 47146 -3132 47382 -2896
rect 51326 707792 51562 708028
rect 51646 707792 51882 708028
rect 51326 707472 51562 707708
rect 51646 707472 51882 707708
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3772 51562 -3536
rect 51646 -3772 51882 -3536
rect 51326 -4092 51562 -3856
rect 51646 -4092 51882 -3856
rect 55826 708752 56062 708988
rect 56146 708752 56382 708988
rect 55826 708432 56062 708668
rect 56146 708432 56382 708668
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4732 56062 -4496
rect 56146 -4732 56382 -4496
rect 55826 -5052 56062 -4816
rect 56146 -5052 56382 -4816
rect 60326 709712 60562 709948
rect 60646 709712 60882 709948
rect 60326 709392 60562 709628
rect 60646 709392 60882 709628
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5692 60562 -5456
rect 60646 -5692 60882 -5456
rect 60326 -6012 60562 -5776
rect 60646 -6012 60882 -5776
rect 64826 710672 65062 710908
rect 65146 710672 65382 710908
rect 64826 710352 65062 710588
rect 65146 710352 65382 710588
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6652 65062 -6416
rect 65146 -6652 65382 -6416
rect 64826 -6972 65062 -6736
rect 65146 -6972 65382 -6736
rect 69326 711632 69562 711868
rect 69646 711632 69882 711868
rect 69326 711312 69562 711548
rect 69646 711312 69882 711548
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7612 69562 -7376
rect 69646 -7612 69882 -7376
rect 69326 -7932 69562 -7696
rect 69646 -7932 69882 -7696
rect 73826 704912 74062 705148
rect 74146 704912 74382 705148
rect 73826 704592 74062 704828
rect 74146 704592 74382 704828
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 705872 78562 706108
rect 78646 705872 78882 706108
rect 78326 705552 78562 705788
rect 78646 705552 78882 705788
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 706832 83062 707068
rect 83146 706832 83382 707068
rect 82826 706512 83062 706748
rect 83146 706512 83382 706748
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 87326 707792 87562 708028
rect 87646 707792 87882 708028
rect 87326 707472 87562 707708
rect 87646 707472 87882 707708
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 91826 708752 92062 708988
rect 92146 708752 92382 708988
rect 91826 708432 92062 708668
rect 92146 708432 92382 708668
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 96326 709712 96562 709948
rect 96646 709712 96882 709948
rect 96326 709392 96562 709628
rect 96646 709392 96882 709628
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 100826 710672 101062 710908
rect 101146 710672 101382 710908
rect 100826 710352 101062 710588
rect 101146 710352 101382 710588
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 105326 711632 105562 711868
rect 105646 711632 105882 711868
rect 105326 711312 105562 711548
rect 105646 711312 105882 711548
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 109826 704912 110062 705148
rect 110146 704912 110382 705148
rect 109826 704592 110062 704828
rect 110146 704592 110382 704828
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 705872 114562 706108
rect 114646 705872 114882 706108
rect 114326 705552 114562 705788
rect 114646 705552 114882 705788
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 706832 119062 707068
rect 119146 706832 119382 707068
rect 118826 706512 119062 706748
rect 119146 706512 119382 706748
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 707792 123562 708028
rect 123646 707792 123882 708028
rect 123326 707472 123562 707708
rect 123646 707472 123882 707708
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -892 74062 -656
rect 74146 -892 74382 -656
rect 73826 -1212 74062 -976
rect 74146 -1212 74382 -976
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1852 78562 -1616
rect 78646 -1852 78882 -1616
rect 78326 -2172 78562 -1936
rect 78646 -2172 78882 -1936
rect 84250 147003 84486 147239
rect 114970 147003 115206 147239
rect 99610 115718 99846 115954
rect 99610 115398 99846 115634
rect 84250 111218 84486 111454
rect 84250 110898 84486 111134
rect 114970 111218 115206 111454
rect 114970 110898 115206 111134
rect 127826 708752 128062 708988
rect 128146 708752 128382 708988
rect 127826 708432 128062 708668
rect 128146 708432 128382 708668
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 82826 -2812 83062 -2576
rect 83146 -2812 83382 -2576
rect 82826 -3132 83062 -2896
rect 83146 -3132 83382 -2896
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 87326 -3772 87562 -3536
rect 87646 -3772 87882 -3536
rect 87326 -4092 87562 -3856
rect 87646 -4092 87882 -3856
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 91826 -4732 92062 -4496
rect 92146 -4732 92382 -4496
rect 91826 -5052 92062 -4816
rect 92146 -5052 92382 -4816
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 96326 -5692 96562 -5456
rect 96646 -5692 96882 -5456
rect 96326 -6012 96562 -5776
rect 96646 -6012 96882 -5776
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 100826 -6652 101062 -6416
rect 101146 -6652 101382 -6416
rect 100826 -6972 101062 -6736
rect 101146 -6972 101382 -6736
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 105326 -7612 105562 -7376
rect 105646 -7612 105882 -7376
rect 105326 -7932 105562 -7696
rect 105646 -7932 105882 -7696
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -892 110062 -656
rect 110146 -892 110382 -656
rect 109826 -1212 110062 -976
rect 110146 -1212 110382 -976
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1852 114562 -1616
rect 114646 -1852 114882 -1616
rect 114326 -2172 114562 -1936
rect 114646 -2172 114882 -1936
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 118826 -2812 119062 -2576
rect 119146 -2812 119382 -2576
rect 118826 -3132 119062 -2896
rect 119146 -3132 119382 -2896
rect 132326 709712 132562 709948
rect 132646 709712 132882 709948
rect 132326 709392 132562 709628
rect 132646 709392 132882 709628
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3772 123562 -3536
rect 123646 -3772 123882 -3536
rect 123326 -4092 123562 -3856
rect 123646 -4092 123882 -3856
rect 127826 -4732 128062 -4496
rect 128146 -4732 128382 -4496
rect 127826 -5052 128062 -4816
rect 128146 -5052 128382 -4816
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5692 132562 -5456
rect 132646 -5692 132882 -5456
rect 132326 -6012 132562 -5776
rect 132646 -6012 132882 -5776
rect 136826 710672 137062 710908
rect 137146 710672 137382 710908
rect 136826 710352 137062 710588
rect 137146 710352 137382 710588
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6652 137062 -6416
rect 137146 -6652 137382 -6416
rect 136826 -6972 137062 -6736
rect 137146 -6972 137382 -6736
rect 141326 711632 141562 711868
rect 141646 711632 141882 711868
rect 141326 711312 141562 711548
rect 141646 711312 141882 711548
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7612 141562 -7376
rect 141646 -7612 141882 -7376
rect 141326 -7932 141562 -7696
rect 141646 -7932 141882 -7696
rect 145826 704912 146062 705148
rect 146146 704912 146382 705148
rect 145826 704592 146062 704828
rect 146146 704592 146382 704828
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -892 146062 -656
rect 146146 -892 146382 -656
rect 145826 -1212 146062 -976
rect 146146 -1212 146382 -976
rect 150326 705872 150562 706108
rect 150646 705872 150882 706108
rect 150326 705552 150562 705788
rect 150646 705552 150882 705788
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1852 150562 -1616
rect 150646 -1852 150882 -1616
rect 150326 -2172 150562 -1936
rect 150646 -2172 150882 -1936
rect 154826 706832 155062 707068
rect 155146 706832 155382 707068
rect 154826 706512 155062 706748
rect 155146 706512 155382 706748
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2812 155062 -2576
rect 155146 -2812 155382 -2576
rect 154826 -3132 155062 -2896
rect 155146 -3132 155382 -2896
rect 159326 707792 159562 708028
rect 159646 707792 159882 708028
rect 159326 707472 159562 707708
rect 159646 707472 159882 707708
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3772 159562 -3536
rect 159646 -3772 159882 -3536
rect 159326 -4092 159562 -3856
rect 159646 -4092 159882 -3856
rect 163826 708752 164062 708988
rect 164146 708752 164382 708988
rect 163826 708432 164062 708668
rect 164146 708432 164382 708668
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4732 164062 -4496
rect 164146 -4732 164382 -4496
rect 163826 -5052 164062 -4816
rect 164146 -5052 164382 -4816
rect 168326 709712 168562 709948
rect 168646 709712 168882 709948
rect 168326 709392 168562 709628
rect 168646 709392 168882 709628
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5692 168562 -5456
rect 168646 -5692 168882 -5456
rect 168326 -6012 168562 -5776
rect 168646 -6012 168882 -5776
rect 172826 710672 173062 710908
rect 173146 710672 173382 710908
rect 172826 710352 173062 710588
rect 173146 710352 173382 710588
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6652 173062 -6416
rect 173146 -6652 173382 -6416
rect 172826 -6972 173062 -6736
rect 173146 -6972 173382 -6736
rect 177326 711632 177562 711868
rect 177646 711632 177882 711868
rect 177326 711312 177562 711548
rect 177646 711312 177882 711548
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7612 177562 -7376
rect 177646 -7612 177882 -7376
rect 177326 -7932 177562 -7696
rect 177646 -7932 177882 -7696
rect 181826 704912 182062 705148
rect 182146 704912 182382 705148
rect 181826 704592 182062 704828
rect 182146 704592 182382 704828
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -892 182062 -656
rect 182146 -892 182382 -656
rect 181826 -1212 182062 -976
rect 182146 -1212 182382 -976
rect 186326 705872 186562 706108
rect 186646 705872 186882 706108
rect 186326 705552 186562 705788
rect 186646 705552 186882 705788
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1852 186562 -1616
rect 186646 -1852 186882 -1616
rect 186326 -2172 186562 -1936
rect 186646 -2172 186882 -1936
rect 190826 706832 191062 707068
rect 191146 706832 191382 707068
rect 190826 706512 191062 706748
rect 191146 706512 191382 706748
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2812 191062 -2576
rect 191146 -2812 191382 -2576
rect 190826 -3132 191062 -2896
rect 191146 -3132 191382 -2896
rect 195326 707792 195562 708028
rect 195646 707792 195882 708028
rect 195326 707472 195562 707708
rect 195646 707472 195882 707708
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3772 195562 -3536
rect 195646 -3772 195882 -3536
rect 195326 -4092 195562 -3856
rect 195646 -4092 195882 -3856
rect 199826 708752 200062 708988
rect 200146 708752 200382 708988
rect 199826 708432 200062 708668
rect 200146 708432 200382 708668
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4732 200062 -4496
rect 200146 -4732 200382 -4496
rect 199826 -5052 200062 -4816
rect 200146 -5052 200382 -4816
rect 204326 709712 204562 709948
rect 204646 709712 204882 709948
rect 204326 709392 204562 709628
rect 204646 709392 204882 709628
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5692 204562 -5456
rect 204646 -5692 204882 -5456
rect 204326 -6012 204562 -5776
rect 204646 -6012 204882 -5776
rect 208826 710672 209062 710908
rect 209146 710672 209382 710908
rect 208826 710352 209062 710588
rect 209146 710352 209382 710588
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6652 209062 -6416
rect 209146 -6652 209382 -6416
rect 208826 -6972 209062 -6736
rect 209146 -6972 209382 -6736
rect 213326 711632 213562 711868
rect 213646 711632 213882 711868
rect 213326 711312 213562 711548
rect 213646 711312 213882 711548
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7612 213562 -7376
rect 213646 -7612 213882 -7376
rect 213326 -7932 213562 -7696
rect 213646 -7932 213882 -7696
rect 217826 704912 218062 705148
rect 218146 704912 218382 705148
rect 217826 704592 218062 704828
rect 218146 704592 218382 704828
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -892 218062 -656
rect 218146 -892 218382 -656
rect 217826 -1212 218062 -976
rect 218146 -1212 218382 -976
rect 222326 705872 222562 706108
rect 222646 705872 222882 706108
rect 222326 705552 222562 705788
rect 222646 705552 222882 705788
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1852 222562 -1616
rect 222646 -1852 222882 -1616
rect 222326 -2172 222562 -1936
rect 222646 -2172 222882 -1936
rect 226826 706832 227062 707068
rect 227146 706832 227382 707068
rect 226826 706512 227062 706748
rect 227146 706512 227382 706748
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2812 227062 -2576
rect 227146 -2812 227382 -2576
rect 226826 -3132 227062 -2896
rect 227146 -3132 227382 -2896
rect 231326 707792 231562 708028
rect 231646 707792 231882 708028
rect 231326 707472 231562 707708
rect 231646 707472 231882 707708
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3772 231562 -3536
rect 231646 -3772 231882 -3536
rect 231326 -4092 231562 -3856
rect 231646 -4092 231882 -3856
rect 235826 708752 236062 708988
rect 236146 708752 236382 708988
rect 235826 708432 236062 708668
rect 236146 708432 236382 708668
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4732 236062 -4496
rect 236146 -4732 236382 -4496
rect 235826 -5052 236062 -4816
rect 236146 -5052 236382 -4816
rect 240326 709712 240562 709948
rect 240646 709712 240882 709948
rect 240326 709392 240562 709628
rect 240646 709392 240882 709628
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5692 240562 -5456
rect 240646 -5692 240882 -5456
rect 240326 -6012 240562 -5776
rect 240646 -6012 240882 -5776
rect 244826 710672 245062 710908
rect 245146 710672 245382 710908
rect 244826 710352 245062 710588
rect 245146 710352 245382 710588
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6652 245062 -6416
rect 245146 -6652 245382 -6416
rect 244826 -6972 245062 -6736
rect 245146 -6972 245382 -6736
rect 249326 711632 249562 711868
rect 249646 711632 249882 711868
rect 249326 711312 249562 711548
rect 249646 711312 249882 711548
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7612 249562 -7376
rect 249646 -7612 249882 -7376
rect 249326 -7932 249562 -7696
rect 249646 -7932 249882 -7696
rect 253826 704912 254062 705148
rect 254146 704912 254382 705148
rect 253826 704592 254062 704828
rect 254146 704592 254382 704828
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -892 254062 -656
rect 254146 -892 254382 -656
rect 253826 -1212 254062 -976
rect 254146 -1212 254382 -976
rect 258326 705872 258562 706108
rect 258646 705872 258882 706108
rect 258326 705552 258562 705788
rect 258646 705552 258882 705788
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1852 258562 -1616
rect 258646 -1852 258882 -1616
rect 258326 -2172 258562 -1936
rect 258646 -2172 258882 -1936
rect 262826 706832 263062 707068
rect 263146 706832 263382 707068
rect 262826 706512 263062 706748
rect 263146 706512 263382 706748
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2812 263062 -2576
rect 263146 -2812 263382 -2576
rect 262826 -3132 263062 -2896
rect 263146 -3132 263382 -2896
rect 267326 707792 267562 708028
rect 267646 707792 267882 708028
rect 267326 707472 267562 707708
rect 267646 707472 267882 707708
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3772 267562 -3536
rect 267646 -3772 267882 -3536
rect 267326 -4092 267562 -3856
rect 267646 -4092 267882 -3856
rect 271826 708752 272062 708988
rect 272146 708752 272382 708988
rect 271826 708432 272062 708668
rect 272146 708432 272382 708668
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4732 272062 -4496
rect 272146 -4732 272382 -4496
rect 271826 -5052 272062 -4816
rect 272146 -5052 272382 -4816
rect 276326 709712 276562 709948
rect 276646 709712 276882 709948
rect 276326 709392 276562 709628
rect 276646 709392 276882 709628
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5692 276562 -5456
rect 276646 -5692 276882 -5456
rect 276326 -6012 276562 -5776
rect 276646 -6012 276882 -5776
rect 280826 710672 281062 710908
rect 281146 710672 281382 710908
rect 280826 710352 281062 710588
rect 281146 710352 281382 710588
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6652 281062 -6416
rect 281146 -6652 281382 -6416
rect 280826 -6972 281062 -6736
rect 281146 -6972 281382 -6736
rect 285326 711632 285562 711868
rect 285646 711632 285882 711868
rect 285326 711312 285562 711548
rect 285646 711312 285882 711548
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7612 285562 -7376
rect 285646 -7612 285882 -7376
rect 285326 -7932 285562 -7696
rect 285646 -7932 285882 -7696
rect 289826 704912 290062 705148
rect 290146 704912 290382 705148
rect 289826 704592 290062 704828
rect 290146 704592 290382 704828
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -892 290062 -656
rect 290146 -892 290382 -656
rect 289826 -1212 290062 -976
rect 290146 -1212 290382 -976
rect 294326 705872 294562 706108
rect 294646 705872 294882 706108
rect 294326 705552 294562 705788
rect 294646 705552 294882 705788
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1852 294562 -1616
rect 294646 -1852 294882 -1616
rect 294326 -2172 294562 -1936
rect 294646 -2172 294882 -1936
rect 298826 706832 299062 707068
rect 299146 706832 299382 707068
rect 298826 706512 299062 706748
rect 299146 706512 299382 706748
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2812 299062 -2576
rect 299146 -2812 299382 -2576
rect 298826 -3132 299062 -2896
rect 299146 -3132 299382 -2896
rect 303326 707792 303562 708028
rect 303646 707792 303882 708028
rect 303326 707472 303562 707708
rect 303646 707472 303882 707708
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3772 303562 -3536
rect 303646 -3772 303882 -3536
rect 303326 -4092 303562 -3856
rect 303646 -4092 303882 -3856
rect 307826 708752 308062 708988
rect 308146 708752 308382 708988
rect 307826 708432 308062 708668
rect 308146 708432 308382 708668
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4732 308062 -4496
rect 308146 -4732 308382 -4496
rect 307826 -5052 308062 -4816
rect 308146 -5052 308382 -4816
rect 312326 709712 312562 709948
rect 312646 709712 312882 709948
rect 312326 709392 312562 709628
rect 312646 709392 312882 709628
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5692 312562 -5456
rect 312646 -5692 312882 -5456
rect 312326 -6012 312562 -5776
rect 312646 -6012 312882 -5776
rect 316826 710672 317062 710908
rect 317146 710672 317382 710908
rect 316826 710352 317062 710588
rect 317146 710352 317382 710588
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6652 317062 -6416
rect 317146 -6652 317382 -6416
rect 316826 -6972 317062 -6736
rect 317146 -6972 317382 -6736
rect 321326 711632 321562 711868
rect 321646 711632 321882 711868
rect 321326 711312 321562 711548
rect 321646 711312 321882 711548
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7612 321562 -7376
rect 321646 -7612 321882 -7376
rect 321326 -7932 321562 -7696
rect 321646 -7932 321882 -7696
rect 325826 704912 326062 705148
rect 326146 704912 326382 705148
rect 325826 704592 326062 704828
rect 326146 704592 326382 704828
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -892 326062 -656
rect 326146 -892 326382 -656
rect 325826 -1212 326062 -976
rect 326146 -1212 326382 -976
rect 330326 705872 330562 706108
rect 330646 705872 330882 706108
rect 330326 705552 330562 705788
rect 330646 705552 330882 705788
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1852 330562 -1616
rect 330646 -1852 330882 -1616
rect 330326 -2172 330562 -1936
rect 330646 -2172 330882 -1936
rect 334826 706832 335062 707068
rect 335146 706832 335382 707068
rect 334826 706512 335062 706748
rect 335146 706512 335382 706748
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2812 335062 -2576
rect 335146 -2812 335382 -2576
rect 334826 -3132 335062 -2896
rect 335146 -3132 335382 -2896
rect 339326 707792 339562 708028
rect 339646 707792 339882 708028
rect 339326 707472 339562 707708
rect 339646 707472 339882 707708
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3772 339562 -3536
rect 339646 -3772 339882 -3536
rect 339326 -4092 339562 -3856
rect 339646 -4092 339882 -3856
rect 343826 708752 344062 708988
rect 344146 708752 344382 708988
rect 343826 708432 344062 708668
rect 344146 708432 344382 708668
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4732 344062 -4496
rect 344146 -4732 344382 -4496
rect 343826 -5052 344062 -4816
rect 344146 -5052 344382 -4816
rect 348326 709712 348562 709948
rect 348646 709712 348882 709948
rect 348326 709392 348562 709628
rect 348646 709392 348882 709628
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5692 348562 -5456
rect 348646 -5692 348882 -5456
rect 348326 -6012 348562 -5776
rect 348646 -6012 348882 -5776
rect 352826 710672 353062 710908
rect 353146 710672 353382 710908
rect 352826 710352 353062 710588
rect 353146 710352 353382 710588
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6652 353062 -6416
rect 353146 -6652 353382 -6416
rect 352826 -6972 353062 -6736
rect 353146 -6972 353382 -6736
rect 357326 711632 357562 711868
rect 357646 711632 357882 711868
rect 357326 711312 357562 711548
rect 357646 711312 357882 711548
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7612 357562 -7376
rect 357646 -7612 357882 -7376
rect 357326 -7932 357562 -7696
rect 357646 -7932 357882 -7696
rect 361826 704912 362062 705148
rect 362146 704912 362382 705148
rect 361826 704592 362062 704828
rect 362146 704592 362382 704828
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -892 362062 -656
rect 362146 -892 362382 -656
rect 361826 -1212 362062 -976
rect 362146 -1212 362382 -976
rect 366326 705872 366562 706108
rect 366646 705872 366882 706108
rect 366326 705552 366562 705788
rect 366646 705552 366882 705788
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1852 366562 -1616
rect 366646 -1852 366882 -1616
rect 366326 -2172 366562 -1936
rect 366646 -2172 366882 -1936
rect 370826 706832 371062 707068
rect 371146 706832 371382 707068
rect 370826 706512 371062 706748
rect 371146 706512 371382 706748
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2812 371062 -2576
rect 371146 -2812 371382 -2576
rect 370826 -3132 371062 -2896
rect 371146 -3132 371382 -2896
rect 375326 707792 375562 708028
rect 375646 707792 375882 708028
rect 375326 707472 375562 707708
rect 375646 707472 375882 707708
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3772 375562 -3536
rect 375646 -3772 375882 -3536
rect 375326 -4092 375562 -3856
rect 375646 -4092 375882 -3856
rect 379826 708752 380062 708988
rect 380146 708752 380382 708988
rect 379826 708432 380062 708668
rect 380146 708432 380382 708668
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4732 380062 -4496
rect 380146 -4732 380382 -4496
rect 379826 -5052 380062 -4816
rect 380146 -5052 380382 -4816
rect 384326 709712 384562 709948
rect 384646 709712 384882 709948
rect 384326 709392 384562 709628
rect 384646 709392 384882 709628
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5692 384562 -5456
rect 384646 -5692 384882 -5456
rect 384326 -6012 384562 -5776
rect 384646 -6012 384882 -5776
rect 388826 710672 389062 710908
rect 389146 710672 389382 710908
rect 388826 710352 389062 710588
rect 389146 710352 389382 710588
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6652 389062 -6416
rect 389146 -6652 389382 -6416
rect 388826 -6972 389062 -6736
rect 389146 -6972 389382 -6736
rect 393326 711632 393562 711868
rect 393646 711632 393882 711868
rect 393326 711312 393562 711548
rect 393646 711312 393882 711548
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7612 393562 -7376
rect 393646 -7612 393882 -7376
rect 393326 -7932 393562 -7696
rect 393646 -7932 393882 -7696
rect 397826 704912 398062 705148
rect 398146 704912 398382 705148
rect 397826 704592 398062 704828
rect 398146 704592 398382 704828
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -892 398062 -656
rect 398146 -892 398382 -656
rect 397826 -1212 398062 -976
rect 398146 -1212 398382 -976
rect 402326 705872 402562 706108
rect 402646 705872 402882 706108
rect 402326 705552 402562 705788
rect 402646 705552 402882 705788
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1852 402562 -1616
rect 402646 -1852 402882 -1616
rect 402326 -2172 402562 -1936
rect 402646 -2172 402882 -1936
rect 406826 706832 407062 707068
rect 407146 706832 407382 707068
rect 406826 706512 407062 706748
rect 407146 706512 407382 706748
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2812 407062 -2576
rect 407146 -2812 407382 -2576
rect 406826 -3132 407062 -2896
rect 407146 -3132 407382 -2896
rect 411326 707792 411562 708028
rect 411646 707792 411882 708028
rect 411326 707472 411562 707708
rect 411646 707472 411882 707708
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3772 411562 -3536
rect 411646 -3772 411882 -3536
rect 411326 -4092 411562 -3856
rect 411646 -4092 411882 -3856
rect 415826 708752 416062 708988
rect 416146 708752 416382 708988
rect 415826 708432 416062 708668
rect 416146 708432 416382 708668
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4732 416062 -4496
rect 416146 -4732 416382 -4496
rect 415826 -5052 416062 -4816
rect 416146 -5052 416382 -4816
rect 420326 709712 420562 709948
rect 420646 709712 420882 709948
rect 420326 709392 420562 709628
rect 420646 709392 420882 709628
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5692 420562 -5456
rect 420646 -5692 420882 -5456
rect 420326 -6012 420562 -5776
rect 420646 -6012 420882 -5776
rect 424826 710672 425062 710908
rect 425146 710672 425382 710908
rect 424826 710352 425062 710588
rect 425146 710352 425382 710588
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6652 425062 -6416
rect 425146 -6652 425382 -6416
rect 424826 -6972 425062 -6736
rect 425146 -6972 425382 -6736
rect 429326 711632 429562 711868
rect 429646 711632 429882 711868
rect 429326 711312 429562 711548
rect 429646 711312 429882 711548
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7612 429562 -7376
rect 429646 -7612 429882 -7376
rect 429326 -7932 429562 -7696
rect 429646 -7932 429882 -7696
rect 433826 704912 434062 705148
rect 434146 704912 434382 705148
rect 433826 704592 434062 704828
rect 434146 704592 434382 704828
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -892 434062 -656
rect 434146 -892 434382 -656
rect 433826 -1212 434062 -976
rect 434146 -1212 434382 -976
rect 438326 705872 438562 706108
rect 438646 705872 438882 706108
rect 438326 705552 438562 705788
rect 438646 705552 438882 705788
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1852 438562 -1616
rect 438646 -1852 438882 -1616
rect 438326 -2172 438562 -1936
rect 438646 -2172 438882 -1936
rect 442826 706832 443062 707068
rect 443146 706832 443382 707068
rect 442826 706512 443062 706748
rect 443146 706512 443382 706748
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2812 443062 -2576
rect 443146 -2812 443382 -2576
rect 442826 -3132 443062 -2896
rect 443146 -3132 443382 -2896
rect 447326 707792 447562 708028
rect 447646 707792 447882 708028
rect 447326 707472 447562 707708
rect 447646 707472 447882 707708
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3772 447562 -3536
rect 447646 -3772 447882 -3536
rect 447326 -4092 447562 -3856
rect 447646 -4092 447882 -3856
rect 451826 708752 452062 708988
rect 452146 708752 452382 708988
rect 451826 708432 452062 708668
rect 452146 708432 452382 708668
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4732 452062 -4496
rect 452146 -4732 452382 -4496
rect 451826 -5052 452062 -4816
rect 452146 -5052 452382 -4816
rect 456326 709712 456562 709948
rect 456646 709712 456882 709948
rect 456326 709392 456562 709628
rect 456646 709392 456882 709628
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5692 456562 -5456
rect 456646 -5692 456882 -5456
rect 456326 -6012 456562 -5776
rect 456646 -6012 456882 -5776
rect 460826 710672 461062 710908
rect 461146 710672 461382 710908
rect 460826 710352 461062 710588
rect 461146 710352 461382 710588
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6652 461062 -6416
rect 461146 -6652 461382 -6416
rect 460826 -6972 461062 -6736
rect 461146 -6972 461382 -6736
rect 465326 711632 465562 711868
rect 465646 711632 465882 711868
rect 465326 711312 465562 711548
rect 465646 711312 465882 711548
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7612 465562 -7376
rect 465646 -7612 465882 -7376
rect 465326 -7932 465562 -7696
rect 465646 -7932 465882 -7696
rect 469826 704912 470062 705148
rect 470146 704912 470382 705148
rect 469826 704592 470062 704828
rect 470146 704592 470382 704828
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -892 470062 -656
rect 470146 -892 470382 -656
rect 469826 -1212 470062 -976
rect 470146 -1212 470382 -976
rect 474326 705872 474562 706108
rect 474646 705872 474882 706108
rect 474326 705552 474562 705788
rect 474646 705552 474882 705788
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1852 474562 -1616
rect 474646 -1852 474882 -1616
rect 474326 -2172 474562 -1936
rect 474646 -2172 474882 -1936
rect 478826 706832 479062 707068
rect 479146 706832 479382 707068
rect 478826 706512 479062 706748
rect 479146 706512 479382 706748
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2812 479062 -2576
rect 479146 -2812 479382 -2576
rect 478826 -3132 479062 -2896
rect 479146 -3132 479382 -2896
rect 483326 707792 483562 708028
rect 483646 707792 483882 708028
rect 483326 707472 483562 707708
rect 483646 707472 483882 707708
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3772 483562 -3536
rect 483646 -3772 483882 -3536
rect 483326 -4092 483562 -3856
rect 483646 -4092 483882 -3856
rect 487826 708752 488062 708988
rect 488146 708752 488382 708988
rect 487826 708432 488062 708668
rect 488146 708432 488382 708668
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4732 488062 -4496
rect 488146 -4732 488382 -4496
rect 487826 -5052 488062 -4816
rect 488146 -5052 488382 -4816
rect 492326 709712 492562 709948
rect 492646 709712 492882 709948
rect 492326 709392 492562 709628
rect 492646 709392 492882 709628
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5692 492562 -5456
rect 492646 -5692 492882 -5456
rect 492326 -6012 492562 -5776
rect 492646 -6012 492882 -5776
rect 496826 710672 497062 710908
rect 497146 710672 497382 710908
rect 496826 710352 497062 710588
rect 497146 710352 497382 710588
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6652 497062 -6416
rect 497146 -6652 497382 -6416
rect 496826 -6972 497062 -6736
rect 497146 -6972 497382 -6736
rect 501326 711632 501562 711868
rect 501646 711632 501882 711868
rect 501326 711312 501562 711548
rect 501646 711312 501882 711548
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7612 501562 -7376
rect 501646 -7612 501882 -7376
rect 501326 -7932 501562 -7696
rect 501646 -7932 501882 -7696
rect 505826 704912 506062 705148
rect 506146 704912 506382 705148
rect 505826 704592 506062 704828
rect 506146 704592 506382 704828
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -892 506062 -656
rect 506146 -892 506382 -656
rect 505826 -1212 506062 -976
rect 506146 -1212 506382 -976
rect 510326 705872 510562 706108
rect 510646 705872 510882 706108
rect 510326 705552 510562 705788
rect 510646 705552 510882 705788
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1852 510562 -1616
rect 510646 -1852 510882 -1616
rect 510326 -2172 510562 -1936
rect 510646 -2172 510882 -1936
rect 514826 706832 515062 707068
rect 515146 706832 515382 707068
rect 514826 706512 515062 706748
rect 515146 706512 515382 706748
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2812 515062 -2576
rect 515146 -2812 515382 -2576
rect 514826 -3132 515062 -2896
rect 515146 -3132 515382 -2896
rect 519326 707792 519562 708028
rect 519646 707792 519882 708028
rect 519326 707472 519562 707708
rect 519646 707472 519882 707708
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3772 519562 -3536
rect 519646 -3772 519882 -3536
rect 519326 -4092 519562 -3856
rect 519646 -4092 519882 -3856
rect 523826 708752 524062 708988
rect 524146 708752 524382 708988
rect 523826 708432 524062 708668
rect 524146 708432 524382 708668
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4732 524062 -4496
rect 524146 -4732 524382 -4496
rect 523826 -5052 524062 -4816
rect 524146 -5052 524382 -4816
rect 528326 709712 528562 709948
rect 528646 709712 528882 709948
rect 528326 709392 528562 709628
rect 528646 709392 528882 709628
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5692 528562 -5456
rect 528646 -5692 528882 -5456
rect 528326 -6012 528562 -5776
rect 528646 -6012 528882 -5776
rect 532826 710672 533062 710908
rect 533146 710672 533382 710908
rect 532826 710352 533062 710588
rect 533146 710352 533382 710588
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6652 533062 -6416
rect 533146 -6652 533382 -6416
rect 532826 -6972 533062 -6736
rect 533146 -6972 533382 -6736
rect 537326 711632 537562 711868
rect 537646 711632 537882 711868
rect 537326 711312 537562 711548
rect 537646 711312 537882 711548
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7612 537562 -7376
rect 537646 -7612 537882 -7376
rect 537326 -7932 537562 -7696
rect 537646 -7932 537882 -7696
rect 541826 704912 542062 705148
rect 542146 704912 542382 705148
rect 541826 704592 542062 704828
rect 542146 704592 542382 704828
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -892 542062 -656
rect 542146 -892 542382 -656
rect 541826 -1212 542062 -976
rect 542146 -1212 542382 -976
rect 546326 705872 546562 706108
rect 546646 705872 546882 706108
rect 546326 705552 546562 705788
rect 546646 705552 546882 705788
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1852 546562 -1616
rect 546646 -1852 546882 -1616
rect 546326 -2172 546562 -1936
rect 546646 -2172 546882 -1936
rect 550826 706832 551062 707068
rect 551146 706832 551382 707068
rect 550826 706512 551062 706748
rect 551146 706512 551382 706748
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2812 551062 -2576
rect 551146 -2812 551382 -2576
rect 550826 -3132 551062 -2896
rect 551146 -3132 551382 -2896
rect 555326 707792 555562 708028
rect 555646 707792 555882 708028
rect 555326 707472 555562 707708
rect 555646 707472 555882 707708
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3772 555562 -3536
rect 555646 -3772 555882 -3536
rect 555326 -4092 555562 -3856
rect 555646 -4092 555882 -3856
rect 559826 708752 560062 708988
rect 560146 708752 560382 708988
rect 559826 708432 560062 708668
rect 560146 708432 560382 708668
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4732 560062 -4496
rect 560146 -4732 560382 -4496
rect 559826 -5052 560062 -4816
rect 560146 -5052 560382 -4816
rect 564326 709712 564562 709948
rect 564646 709712 564882 709948
rect 564326 709392 564562 709628
rect 564646 709392 564882 709628
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5692 564562 -5456
rect 564646 -5692 564882 -5456
rect 564326 -6012 564562 -5776
rect 564646 -6012 564882 -5776
rect 568826 710672 569062 710908
rect 569146 710672 569382 710908
rect 568826 710352 569062 710588
rect 569146 710352 569382 710588
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6652 569062 -6416
rect 569146 -6652 569382 -6416
rect 568826 -6972 569062 -6736
rect 569146 -6972 569382 -6736
rect 573326 711632 573562 711868
rect 573646 711632 573882 711868
rect 573326 711312 573562 711548
rect 573646 711312 573882 711548
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7612 573562 -7376
rect 573646 -7612 573882 -7376
rect 573326 -7932 573562 -7696
rect 573646 -7932 573882 -7696
rect 577826 704912 578062 705148
rect 578146 704912 578382 705148
rect 577826 704592 578062 704828
rect 578146 704592 578382 704828
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -892 578062 -656
rect 578146 -892 578382 -656
rect 577826 -1212 578062 -976
rect 578146 -1212 578382 -976
rect 592372 711632 592608 711868
rect 592692 711632 592928 711868
rect 592372 711312 592608 711548
rect 592692 711312 592928 711548
rect 591412 710672 591648 710908
rect 591732 710672 591968 710908
rect 591412 710352 591648 710588
rect 591732 710352 591968 710588
rect 590452 709712 590688 709948
rect 590772 709712 591008 709948
rect 590452 709392 590688 709628
rect 590772 709392 591008 709628
rect 589492 708752 589728 708988
rect 589812 708752 590048 708988
rect 589492 708432 589728 708668
rect 589812 708432 590048 708668
rect 588532 707792 588768 708028
rect 588852 707792 589088 708028
rect 588532 707472 588768 707708
rect 588852 707472 589088 707708
rect 587572 706832 587808 707068
rect 587892 706832 588128 707068
rect 587572 706512 587808 706748
rect 587892 706512 588128 706748
rect 582326 705872 582562 706108
rect 582646 705872 582882 706108
rect 582326 705552 582562 705788
rect 582646 705552 582882 705788
rect 586612 705872 586848 706108
rect 586932 705872 587168 706108
rect 586612 705552 586848 705788
rect 586932 705552 587168 705788
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585652 704912 585888 705148
rect 585972 704912 586208 705148
rect 585652 704592 585888 704828
rect 585972 704592 586208 704828
rect 585652 687218 585888 687454
rect 585972 687218 586208 687454
rect 585652 686898 585888 687134
rect 585972 686898 586208 687134
rect 585652 651218 585888 651454
rect 585972 651218 586208 651454
rect 585652 650898 585888 651134
rect 585972 650898 586208 651134
rect 585652 615218 585888 615454
rect 585972 615218 586208 615454
rect 585652 614898 585888 615134
rect 585972 614898 586208 615134
rect 585652 579218 585888 579454
rect 585972 579218 586208 579454
rect 585652 578898 585888 579134
rect 585972 578898 586208 579134
rect 585652 543218 585888 543454
rect 585972 543218 586208 543454
rect 585652 542898 585888 543134
rect 585972 542898 586208 543134
rect 585652 507218 585888 507454
rect 585972 507218 586208 507454
rect 585652 506898 585888 507134
rect 585972 506898 586208 507134
rect 585652 471218 585888 471454
rect 585972 471218 586208 471454
rect 585652 470898 585888 471134
rect 585972 470898 586208 471134
rect 585652 435218 585888 435454
rect 585972 435218 586208 435454
rect 585652 434898 585888 435134
rect 585972 434898 586208 435134
rect 585652 399218 585888 399454
rect 585972 399218 586208 399454
rect 585652 398898 585888 399134
rect 585972 398898 586208 399134
rect 585652 363218 585888 363454
rect 585972 363218 586208 363454
rect 585652 362898 585888 363134
rect 585972 362898 586208 363134
rect 585652 327218 585888 327454
rect 585972 327218 586208 327454
rect 585652 326898 585888 327134
rect 585972 326898 586208 327134
rect 585652 291218 585888 291454
rect 585972 291218 586208 291454
rect 585652 290898 585888 291134
rect 585972 290898 586208 291134
rect 585652 255218 585888 255454
rect 585972 255218 586208 255454
rect 585652 254898 585888 255134
rect 585972 254898 586208 255134
rect 585652 219218 585888 219454
rect 585972 219218 586208 219454
rect 585652 218898 585888 219134
rect 585972 218898 586208 219134
rect 585652 183218 585888 183454
rect 585972 183218 586208 183454
rect 585652 182898 585888 183134
rect 585972 182898 586208 183134
rect 585652 147218 585888 147454
rect 585972 147218 586208 147454
rect 585652 146898 585888 147134
rect 585972 146898 586208 147134
rect 585652 111218 585888 111454
rect 585972 111218 586208 111454
rect 585652 110898 585888 111134
rect 585972 110898 586208 111134
rect 585652 75218 585888 75454
rect 585972 75218 586208 75454
rect 585652 74898 585888 75134
rect 585972 74898 586208 75134
rect 585652 39218 585888 39454
rect 585972 39218 586208 39454
rect 585652 38898 585888 39134
rect 585972 38898 586208 39134
rect 585652 3218 585888 3454
rect 585972 3218 586208 3454
rect 585652 2898 585888 3134
rect 585972 2898 586208 3134
rect 585652 -892 585888 -656
rect 585972 -892 586208 -656
rect 585652 -1212 585888 -976
rect 585972 -1212 586208 -976
rect 586612 691718 586848 691954
rect 586932 691718 587168 691954
rect 586612 691398 586848 691634
rect 586932 691398 587168 691634
rect 586612 655718 586848 655954
rect 586932 655718 587168 655954
rect 586612 655398 586848 655634
rect 586932 655398 587168 655634
rect 586612 619718 586848 619954
rect 586932 619718 587168 619954
rect 586612 619398 586848 619634
rect 586932 619398 587168 619634
rect 586612 583718 586848 583954
rect 586932 583718 587168 583954
rect 586612 583398 586848 583634
rect 586932 583398 587168 583634
rect 586612 547718 586848 547954
rect 586932 547718 587168 547954
rect 586612 547398 586848 547634
rect 586932 547398 587168 547634
rect 586612 511718 586848 511954
rect 586932 511718 587168 511954
rect 586612 511398 586848 511634
rect 586932 511398 587168 511634
rect 586612 475718 586848 475954
rect 586932 475718 587168 475954
rect 586612 475398 586848 475634
rect 586932 475398 587168 475634
rect 586612 439718 586848 439954
rect 586932 439718 587168 439954
rect 586612 439398 586848 439634
rect 586932 439398 587168 439634
rect 586612 403718 586848 403954
rect 586932 403718 587168 403954
rect 586612 403398 586848 403634
rect 586932 403398 587168 403634
rect 586612 367718 586848 367954
rect 586932 367718 587168 367954
rect 586612 367398 586848 367634
rect 586932 367398 587168 367634
rect 586612 331718 586848 331954
rect 586932 331718 587168 331954
rect 586612 331398 586848 331634
rect 586932 331398 587168 331634
rect 586612 295718 586848 295954
rect 586932 295718 587168 295954
rect 586612 295398 586848 295634
rect 586932 295398 587168 295634
rect 586612 259718 586848 259954
rect 586932 259718 587168 259954
rect 586612 259398 586848 259634
rect 586932 259398 587168 259634
rect 586612 223718 586848 223954
rect 586932 223718 587168 223954
rect 586612 223398 586848 223634
rect 586932 223398 587168 223634
rect 586612 187718 586848 187954
rect 586932 187718 587168 187954
rect 586612 187398 586848 187634
rect 586932 187398 587168 187634
rect 586612 151718 586848 151954
rect 586932 151718 587168 151954
rect 586612 151398 586848 151634
rect 586932 151398 587168 151634
rect 586612 115718 586848 115954
rect 586932 115718 587168 115954
rect 586612 115398 586848 115634
rect 586932 115398 587168 115634
rect 586612 79718 586848 79954
rect 586932 79718 587168 79954
rect 586612 79398 586848 79634
rect 586932 79398 587168 79634
rect 586612 43718 586848 43954
rect 586932 43718 587168 43954
rect 586612 43398 586848 43634
rect 586932 43398 587168 43634
rect 586612 7718 586848 7954
rect 586932 7718 587168 7954
rect 586612 7398 586848 7634
rect 586932 7398 587168 7634
rect 582326 -1852 582562 -1616
rect 582646 -1852 582882 -1616
rect 582326 -2172 582562 -1936
rect 582646 -2172 582882 -1936
rect 586612 -1852 586848 -1616
rect 586932 -1852 587168 -1616
rect 586612 -2172 586848 -1936
rect 586932 -2172 587168 -1936
rect 587572 696218 587808 696454
rect 587892 696218 588128 696454
rect 587572 695898 587808 696134
rect 587892 695898 588128 696134
rect 587572 660218 587808 660454
rect 587892 660218 588128 660454
rect 587572 659898 587808 660134
rect 587892 659898 588128 660134
rect 587572 624218 587808 624454
rect 587892 624218 588128 624454
rect 587572 623898 587808 624134
rect 587892 623898 588128 624134
rect 587572 588218 587808 588454
rect 587892 588218 588128 588454
rect 587572 587898 587808 588134
rect 587892 587898 588128 588134
rect 587572 552218 587808 552454
rect 587892 552218 588128 552454
rect 587572 551898 587808 552134
rect 587892 551898 588128 552134
rect 587572 516218 587808 516454
rect 587892 516218 588128 516454
rect 587572 515898 587808 516134
rect 587892 515898 588128 516134
rect 587572 480218 587808 480454
rect 587892 480218 588128 480454
rect 587572 479898 587808 480134
rect 587892 479898 588128 480134
rect 587572 444218 587808 444454
rect 587892 444218 588128 444454
rect 587572 443898 587808 444134
rect 587892 443898 588128 444134
rect 587572 408218 587808 408454
rect 587892 408218 588128 408454
rect 587572 407898 587808 408134
rect 587892 407898 588128 408134
rect 587572 372218 587808 372454
rect 587892 372218 588128 372454
rect 587572 371898 587808 372134
rect 587892 371898 588128 372134
rect 587572 336218 587808 336454
rect 587892 336218 588128 336454
rect 587572 335898 587808 336134
rect 587892 335898 588128 336134
rect 587572 300218 587808 300454
rect 587892 300218 588128 300454
rect 587572 299898 587808 300134
rect 587892 299898 588128 300134
rect 587572 264218 587808 264454
rect 587892 264218 588128 264454
rect 587572 263898 587808 264134
rect 587892 263898 588128 264134
rect 587572 228218 587808 228454
rect 587892 228218 588128 228454
rect 587572 227898 587808 228134
rect 587892 227898 588128 228134
rect 587572 192218 587808 192454
rect 587892 192218 588128 192454
rect 587572 191898 587808 192134
rect 587892 191898 588128 192134
rect 587572 156218 587808 156454
rect 587892 156218 588128 156454
rect 587572 155898 587808 156134
rect 587892 155898 588128 156134
rect 587572 120218 587808 120454
rect 587892 120218 588128 120454
rect 587572 119898 587808 120134
rect 587892 119898 588128 120134
rect 587572 84218 587808 84454
rect 587892 84218 588128 84454
rect 587572 83898 587808 84134
rect 587892 83898 588128 84134
rect 587572 48218 587808 48454
rect 587892 48218 588128 48454
rect 587572 47898 587808 48134
rect 587892 47898 588128 48134
rect 587572 12218 587808 12454
rect 587892 12218 588128 12454
rect 587572 11898 587808 12134
rect 587892 11898 588128 12134
rect 587572 -2812 587808 -2576
rect 587892 -2812 588128 -2576
rect 587572 -3132 587808 -2896
rect 587892 -3132 588128 -2896
rect 588532 700718 588768 700954
rect 588852 700718 589088 700954
rect 588532 700398 588768 700634
rect 588852 700398 589088 700634
rect 588532 664718 588768 664954
rect 588852 664718 589088 664954
rect 588532 664398 588768 664634
rect 588852 664398 589088 664634
rect 588532 628718 588768 628954
rect 588852 628718 589088 628954
rect 588532 628398 588768 628634
rect 588852 628398 589088 628634
rect 588532 592718 588768 592954
rect 588852 592718 589088 592954
rect 588532 592398 588768 592634
rect 588852 592398 589088 592634
rect 588532 556718 588768 556954
rect 588852 556718 589088 556954
rect 588532 556398 588768 556634
rect 588852 556398 589088 556634
rect 588532 520718 588768 520954
rect 588852 520718 589088 520954
rect 588532 520398 588768 520634
rect 588852 520398 589088 520634
rect 588532 484718 588768 484954
rect 588852 484718 589088 484954
rect 588532 484398 588768 484634
rect 588852 484398 589088 484634
rect 588532 448718 588768 448954
rect 588852 448718 589088 448954
rect 588532 448398 588768 448634
rect 588852 448398 589088 448634
rect 588532 412718 588768 412954
rect 588852 412718 589088 412954
rect 588532 412398 588768 412634
rect 588852 412398 589088 412634
rect 588532 376718 588768 376954
rect 588852 376718 589088 376954
rect 588532 376398 588768 376634
rect 588852 376398 589088 376634
rect 588532 340718 588768 340954
rect 588852 340718 589088 340954
rect 588532 340398 588768 340634
rect 588852 340398 589088 340634
rect 588532 304718 588768 304954
rect 588852 304718 589088 304954
rect 588532 304398 588768 304634
rect 588852 304398 589088 304634
rect 588532 268718 588768 268954
rect 588852 268718 589088 268954
rect 588532 268398 588768 268634
rect 588852 268398 589088 268634
rect 588532 232718 588768 232954
rect 588852 232718 589088 232954
rect 588532 232398 588768 232634
rect 588852 232398 589088 232634
rect 588532 196718 588768 196954
rect 588852 196718 589088 196954
rect 588532 196398 588768 196634
rect 588852 196398 589088 196634
rect 588532 160718 588768 160954
rect 588852 160718 589088 160954
rect 588532 160398 588768 160634
rect 588852 160398 589088 160634
rect 588532 124718 588768 124954
rect 588852 124718 589088 124954
rect 588532 124398 588768 124634
rect 588852 124398 589088 124634
rect 588532 88718 588768 88954
rect 588852 88718 589088 88954
rect 588532 88398 588768 88634
rect 588852 88398 589088 88634
rect 588532 52718 588768 52954
rect 588852 52718 589088 52954
rect 588532 52398 588768 52634
rect 588852 52398 589088 52634
rect 588532 16718 588768 16954
rect 588852 16718 589088 16954
rect 588532 16398 588768 16634
rect 588852 16398 589088 16634
rect 588532 -3772 588768 -3536
rect 588852 -3772 589088 -3536
rect 588532 -4092 588768 -3856
rect 588852 -4092 589088 -3856
rect 589492 669218 589728 669454
rect 589812 669218 590048 669454
rect 589492 668898 589728 669134
rect 589812 668898 590048 669134
rect 589492 633218 589728 633454
rect 589812 633218 590048 633454
rect 589492 632898 589728 633134
rect 589812 632898 590048 633134
rect 589492 597218 589728 597454
rect 589812 597218 590048 597454
rect 589492 596898 589728 597134
rect 589812 596898 590048 597134
rect 589492 561218 589728 561454
rect 589812 561218 590048 561454
rect 589492 560898 589728 561134
rect 589812 560898 590048 561134
rect 589492 525218 589728 525454
rect 589812 525218 590048 525454
rect 589492 524898 589728 525134
rect 589812 524898 590048 525134
rect 589492 489218 589728 489454
rect 589812 489218 590048 489454
rect 589492 488898 589728 489134
rect 589812 488898 590048 489134
rect 589492 453218 589728 453454
rect 589812 453218 590048 453454
rect 589492 452898 589728 453134
rect 589812 452898 590048 453134
rect 589492 417218 589728 417454
rect 589812 417218 590048 417454
rect 589492 416898 589728 417134
rect 589812 416898 590048 417134
rect 589492 381218 589728 381454
rect 589812 381218 590048 381454
rect 589492 380898 589728 381134
rect 589812 380898 590048 381134
rect 589492 345218 589728 345454
rect 589812 345218 590048 345454
rect 589492 344898 589728 345134
rect 589812 344898 590048 345134
rect 589492 309218 589728 309454
rect 589812 309218 590048 309454
rect 589492 308898 589728 309134
rect 589812 308898 590048 309134
rect 589492 273218 589728 273454
rect 589812 273218 590048 273454
rect 589492 272898 589728 273134
rect 589812 272898 590048 273134
rect 589492 237218 589728 237454
rect 589812 237218 590048 237454
rect 589492 236898 589728 237134
rect 589812 236898 590048 237134
rect 589492 201218 589728 201454
rect 589812 201218 590048 201454
rect 589492 200898 589728 201134
rect 589812 200898 590048 201134
rect 589492 165218 589728 165454
rect 589812 165218 590048 165454
rect 589492 164898 589728 165134
rect 589812 164898 590048 165134
rect 589492 129218 589728 129454
rect 589812 129218 590048 129454
rect 589492 128898 589728 129134
rect 589812 128898 590048 129134
rect 589492 93218 589728 93454
rect 589812 93218 590048 93454
rect 589492 92898 589728 93134
rect 589812 92898 590048 93134
rect 589492 57218 589728 57454
rect 589812 57218 590048 57454
rect 589492 56898 589728 57134
rect 589812 56898 590048 57134
rect 589492 21218 589728 21454
rect 589812 21218 590048 21454
rect 589492 20898 589728 21134
rect 589812 20898 590048 21134
rect 589492 -4732 589728 -4496
rect 589812 -4732 590048 -4496
rect 589492 -5052 589728 -4816
rect 589812 -5052 590048 -4816
rect 590452 673718 590688 673954
rect 590772 673718 591008 673954
rect 590452 673398 590688 673634
rect 590772 673398 591008 673634
rect 590452 637718 590688 637954
rect 590772 637718 591008 637954
rect 590452 637398 590688 637634
rect 590772 637398 591008 637634
rect 590452 601718 590688 601954
rect 590772 601718 591008 601954
rect 590452 601398 590688 601634
rect 590772 601398 591008 601634
rect 590452 565718 590688 565954
rect 590772 565718 591008 565954
rect 590452 565398 590688 565634
rect 590772 565398 591008 565634
rect 590452 529718 590688 529954
rect 590772 529718 591008 529954
rect 590452 529398 590688 529634
rect 590772 529398 591008 529634
rect 590452 493718 590688 493954
rect 590772 493718 591008 493954
rect 590452 493398 590688 493634
rect 590772 493398 591008 493634
rect 590452 457718 590688 457954
rect 590772 457718 591008 457954
rect 590452 457398 590688 457634
rect 590772 457398 591008 457634
rect 590452 421718 590688 421954
rect 590772 421718 591008 421954
rect 590452 421398 590688 421634
rect 590772 421398 591008 421634
rect 590452 385718 590688 385954
rect 590772 385718 591008 385954
rect 590452 385398 590688 385634
rect 590772 385398 591008 385634
rect 590452 349718 590688 349954
rect 590772 349718 591008 349954
rect 590452 349398 590688 349634
rect 590772 349398 591008 349634
rect 590452 313718 590688 313954
rect 590772 313718 591008 313954
rect 590452 313398 590688 313634
rect 590772 313398 591008 313634
rect 590452 277718 590688 277954
rect 590772 277718 591008 277954
rect 590452 277398 590688 277634
rect 590772 277398 591008 277634
rect 590452 241718 590688 241954
rect 590772 241718 591008 241954
rect 590452 241398 590688 241634
rect 590772 241398 591008 241634
rect 590452 205718 590688 205954
rect 590772 205718 591008 205954
rect 590452 205398 590688 205634
rect 590772 205398 591008 205634
rect 590452 169718 590688 169954
rect 590772 169718 591008 169954
rect 590452 169398 590688 169634
rect 590772 169398 591008 169634
rect 590452 133718 590688 133954
rect 590772 133718 591008 133954
rect 590452 133398 590688 133634
rect 590772 133398 591008 133634
rect 590452 97718 590688 97954
rect 590772 97718 591008 97954
rect 590452 97398 590688 97634
rect 590772 97398 591008 97634
rect 590452 61718 590688 61954
rect 590772 61718 591008 61954
rect 590452 61398 590688 61634
rect 590772 61398 591008 61634
rect 590452 25718 590688 25954
rect 590772 25718 591008 25954
rect 590452 25398 590688 25634
rect 590772 25398 591008 25634
rect 590452 -5692 590688 -5456
rect 590772 -5692 591008 -5456
rect 590452 -6012 590688 -5776
rect 590772 -6012 591008 -5776
rect 591412 678218 591648 678454
rect 591732 678218 591968 678454
rect 591412 677898 591648 678134
rect 591732 677898 591968 678134
rect 591412 642218 591648 642454
rect 591732 642218 591968 642454
rect 591412 641898 591648 642134
rect 591732 641898 591968 642134
rect 591412 606218 591648 606454
rect 591732 606218 591968 606454
rect 591412 605898 591648 606134
rect 591732 605898 591968 606134
rect 591412 570218 591648 570454
rect 591732 570218 591968 570454
rect 591412 569898 591648 570134
rect 591732 569898 591968 570134
rect 591412 534218 591648 534454
rect 591732 534218 591968 534454
rect 591412 533898 591648 534134
rect 591732 533898 591968 534134
rect 591412 498218 591648 498454
rect 591732 498218 591968 498454
rect 591412 497898 591648 498134
rect 591732 497898 591968 498134
rect 591412 462218 591648 462454
rect 591732 462218 591968 462454
rect 591412 461898 591648 462134
rect 591732 461898 591968 462134
rect 591412 426218 591648 426454
rect 591732 426218 591968 426454
rect 591412 425898 591648 426134
rect 591732 425898 591968 426134
rect 591412 390218 591648 390454
rect 591732 390218 591968 390454
rect 591412 389898 591648 390134
rect 591732 389898 591968 390134
rect 591412 354218 591648 354454
rect 591732 354218 591968 354454
rect 591412 353898 591648 354134
rect 591732 353898 591968 354134
rect 591412 318218 591648 318454
rect 591732 318218 591968 318454
rect 591412 317898 591648 318134
rect 591732 317898 591968 318134
rect 591412 282218 591648 282454
rect 591732 282218 591968 282454
rect 591412 281898 591648 282134
rect 591732 281898 591968 282134
rect 591412 246218 591648 246454
rect 591732 246218 591968 246454
rect 591412 245898 591648 246134
rect 591732 245898 591968 246134
rect 591412 210218 591648 210454
rect 591732 210218 591968 210454
rect 591412 209898 591648 210134
rect 591732 209898 591968 210134
rect 591412 174218 591648 174454
rect 591732 174218 591968 174454
rect 591412 173898 591648 174134
rect 591732 173898 591968 174134
rect 591412 138218 591648 138454
rect 591732 138218 591968 138454
rect 591412 137898 591648 138134
rect 591732 137898 591968 138134
rect 591412 102218 591648 102454
rect 591732 102218 591968 102454
rect 591412 101898 591648 102134
rect 591732 101898 591968 102134
rect 591412 66218 591648 66454
rect 591732 66218 591968 66454
rect 591412 65898 591648 66134
rect 591732 65898 591968 66134
rect 591412 30218 591648 30454
rect 591732 30218 591968 30454
rect 591412 29898 591648 30134
rect 591732 29898 591968 30134
rect 591412 -6652 591648 -6416
rect 591732 -6652 591968 -6416
rect 591412 -6972 591648 -6736
rect 591732 -6972 591968 -6736
rect 592372 682718 592608 682954
rect 592692 682718 592928 682954
rect 592372 682398 592608 682634
rect 592692 682398 592928 682634
rect 592372 646718 592608 646954
rect 592692 646718 592928 646954
rect 592372 646398 592608 646634
rect 592692 646398 592928 646634
rect 592372 610718 592608 610954
rect 592692 610718 592928 610954
rect 592372 610398 592608 610634
rect 592692 610398 592928 610634
rect 592372 574718 592608 574954
rect 592692 574718 592928 574954
rect 592372 574398 592608 574634
rect 592692 574398 592928 574634
rect 592372 538718 592608 538954
rect 592692 538718 592928 538954
rect 592372 538398 592608 538634
rect 592692 538398 592928 538634
rect 592372 502718 592608 502954
rect 592692 502718 592928 502954
rect 592372 502398 592608 502634
rect 592692 502398 592928 502634
rect 592372 466718 592608 466954
rect 592692 466718 592928 466954
rect 592372 466398 592608 466634
rect 592692 466398 592928 466634
rect 592372 430718 592608 430954
rect 592692 430718 592928 430954
rect 592372 430398 592608 430634
rect 592692 430398 592928 430634
rect 592372 394718 592608 394954
rect 592692 394718 592928 394954
rect 592372 394398 592608 394634
rect 592692 394398 592928 394634
rect 592372 358718 592608 358954
rect 592692 358718 592928 358954
rect 592372 358398 592608 358634
rect 592692 358398 592928 358634
rect 592372 322718 592608 322954
rect 592692 322718 592928 322954
rect 592372 322398 592608 322634
rect 592692 322398 592928 322634
rect 592372 286718 592608 286954
rect 592692 286718 592928 286954
rect 592372 286398 592608 286634
rect 592692 286398 592928 286634
rect 592372 250718 592608 250954
rect 592692 250718 592928 250954
rect 592372 250398 592608 250634
rect 592692 250398 592928 250634
rect 592372 214718 592608 214954
rect 592692 214718 592928 214954
rect 592372 214398 592608 214634
rect 592692 214398 592928 214634
rect 592372 178718 592608 178954
rect 592692 178718 592928 178954
rect 592372 178398 592608 178634
rect 592692 178398 592928 178634
rect 592372 142718 592608 142954
rect 592692 142718 592928 142954
rect 592372 142398 592608 142634
rect 592692 142398 592928 142634
rect 592372 106718 592608 106954
rect 592692 106718 592928 106954
rect 592372 106398 592608 106634
rect 592692 106398 592928 106634
rect 592372 70718 592608 70954
rect 592692 70718 592928 70954
rect 592372 70398 592608 70634
rect 592692 70398 592928 70634
rect 592372 34718 592608 34954
rect 592692 34718 592928 34954
rect 592372 34398 592608 34634
rect 592692 34398 592928 34634
rect 592372 -7612 592608 -7376
rect 592692 -7612 592928 -7376
rect 592372 -7932 592608 -7696
rect 592692 -7932 592928 -7696
<< metal5 >>
rect -9036 711868 592960 711900
rect -9036 711632 -9004 711868
rect -8768 711632 -8684 711868
rect -8448 711632 33326 711868
rect 33562 711632 33646 711868
rect 33882 711632 69326 711868
rect 69562 711632 69646 711868
rect 69882 711632 105326 711868
rect 105562 711632 105646 711868
rect 105882 711632 141326 711868
rect 141562 711632 141646 711868
rect 141882 711632 177326 711868
rect 177562 711632 177646 711868
rect 177882 711632 213326 711868
rect 213562 711632 213646 711868
rect 213882 711632 249326 711868
rect 249562 711632 249646 711868
rect 249882 711632 285326 711868
rect 285562 711632 285646 711868
rect 285882 711632 321326 711868
rect 321562 711632 321646 711868
rect 321882 711632 357326 711868
rect 357562 711632 357646 711868
rect 357882 711632 393326 711868
rect 393562 711632 393646 711868
rect 393882 711632 429326 711868
rect 429562 711632 429646 711868
rect 429882 711632 465326 711868
rect 465562 711632 465646 711868
rect 465882 711632 501326 711868
rect 501562 711632 501646 711868
rect 501882 711632 537326 711868
rect 537562 711632 537646 711868
rect 537882 711632 573326 711868
rect 573562 711632 573646 711868
rect 573882 711632 592372 711868
rect 592608 711632 592692 711868
rect 592928 711632 592960 711868
rect -9036 711548 592960 711632
rect -9036 711312 -9004 711548
rect -8768 711312 -8684 711548
rect -8448 711312 33326 711548
rect 33562 711312 33646 711548
rect 33882 711312 69326 711548
rect 69562 711312 69646 711548
rect 69882 711312 105326 711548
rect 105562 711312 105646 711548
rect 105882 711312 141326 711548
rect 141562 711312 141646 711548
rect 141882 711312 177326 711548
rect 177562 711312 177646 711548
rect 177882 711312 213326 711548
rect 213562 711312 213646 711548
rect 213882 711312 249326 711548
rect 249562 711312 249646 711548
rect 249882 711312 285326 711548
rect 285562 711312 285646 711548
rect 285882 711312 321326 711548
rect 321562 711312 321646 711548
rect 321882 711312 357326 711548
rect 357562 711312 357646 711548
rect 357882 711312 393326 711548
rect 393562 711312 393646 711548
rect 393882 711312 429326 711548
rect 429562 711312 429646 711548
rect 429882 711312 465326 711548
rect 465562 711312 465646 711548
rect 465882 711312 501326 711548
rect 501562 711312 501646 711548
rect 501882 711312 537326 711548
rect 537562 711312 537646 711548
rect 537882 711312 573326 711548
rect 573562 711312 573646 711548
rect 573882 711312 592372 711548
rect 592608 711312 592692 711548
rect 592928 711312 592960 711548
rect -9036 711280 592960 711312
rect -8076 710908 592000 710940
rect -8076 710672 -8044 710908
rect -7808 710672 -7724 710908
rect -7488 710672 28826 710908
rect 29062 710672 29146 710908
rect 29382 710672 64826 710908
rect 65062 710672 65146 710908
rect 65382 710672 100826 710908
rect 101062 710672 101146 710908
rect 101382 710672 136826 710908
rect 137062 710672 137146 710908
rect 137382 710672 172826 710908
rect 173062 710672 173146 710908
rect 173382 710672 208826 710908
rect 209062 710672 209146 710908
rect 209382 710672 244826 710908
rect 245062 710672 245146 710908
rect 245382 710672 280826 710908
rect 281062 710672 281146 710908
rect 281382 710672 316826 710908
rect 317062 710672 317146 710908
rect 317382 710672 352826 710908
rect 353062 710672 353146 710908
rect 353382 710672 388826 710908
rect 389062 710672 389146 710908
rect 389382 710672 424826 710908
rect 425062 710672 425146 710908
rect 425382 710672 460826 710908
rect 461062 710672 461146 710908
rect 461382 710672 496826 710908
rect 497062 710672 497146 710908
rect 497382 710672 532826 710908
rect 533062 710672 533146 710908
rect 533382 710672 568826 710908
rect 569062 710672 569146 710908
rect 569382 710672 591412 710908
rect 591648 710672 591732 710908
rect 591968 710672 592000 710908
rect -8076 710588 592000 710672
rect -8076 710352 -8044 710588
rect -7808 710352 -7724 710588
rect -7488 710352 28826 710588
rect 29062 710352 29146 710588
rect 29382 710352 64826 710588
rect 65062 710352 65146 710588
rect 65382 710352 100826 710588
rect 101062 710352 101146 710588
rect 101382 710352 136826 710588
rect 137062 710352 137146 710588
rect 137382 710352 172826 710588
rect 173062 710352 173146 710588
rect 173382 710352 208826 710588
rect 209062 710352 209146 710588
rect 209382 710352 244826 710588
rect 245062 710352 245146 710588
rect 245382 710352 280826 710588
rect 281062 710352 281146 710588
rect 281382 710352 316826 710588
rect 317062 710352 317146 710588
rect 317382 710352 352826 710588
rect 353062 710352 353146 710588
rect 353382 710352 388826 710588
rect 389062 710352 389146 710588
rect 389382 710352 424826 710588
rect 425062 710352 425146 710588
rect 425382 710352 460826 710588
rect 461062 710352 461146 710588
rect 461382 710352 496826 710588
rect 497062 710352 497146 710588
rect 497382 710352 532826 710588
rect 533062 710352 533146 710588
rect 533382 710352 568826 710588
rect 569062 710352 569146 710588
rect 569382 710352 591412 710588
rect 591648 710352 591732 710588
rect 591968 710352 592000 710588
rect -8076 710320 592000 710352
rect -7116 709948 591040 709980
rect -7116 709712 -7084 709948
rect -6848 709712 -6764 709948
rect -6528 709712 24326 709948
rect 24562 709712 24646 709948
rect 24882 709712 60326 709948
rect 60562 709712 60646 709948
rect 60882 709712 96326 709948
rect 96562 709712 96646 709948
rect 96882 709712 132326 709948
rect 132562 709712 132646 709948
rect 132882 709712 168326 709948
rect 168562 709712 168646 709948
rect 168882 709712 204326 709948
rect 204562 709712 204646 709948
rect 204882 709712 240326 709948
rect 240562 709712 240646 709948
rect 240882 709712 276326 709948
rect 276562 709712 276646 709948
rect 276882 709712 312326 709948
rect 312562 709712 312646 709948
rect 312882 709712 348326 709948
rect 348562 709712 348646 709948
rect 348882 709712 384326 709948
rect 384562 709712 384646 709948
rect 384882 709712 420326 709948
rect 420562 709712 420646 709948
rect 420882 709712 456326 709948
rect 456562 709712 456646 709948
rect 456882 709712 492326 709948
rect 492562 709712 492646 709948
rect 492882 709712 528326 709948
rect 528562 709712 528646 709948
rect 528882 709712 564326 709948
rect 564562 709712 564646 709948
rect 564882 709712 590452 709948
rect 590688 709712 590772 709948
rect 591008 709712 591040 709948
rect -7116 709628 591040 709712
rect -7116 709392 -7084 709628
rect -6848 709392 -6764 709628
rect -6528 709392 24326 709628
rect 24562 709392 24646 709628
rect 24882 709392 60326 709628
rect 60562 709392 60646 709628
rect 60882 709392 96326 709628
rect 96562 709392 96646 709628
rect 96882 709392 132326 709628
rect 132562 709392 132646 709628
rect 132882 709392 168326 709628
rect 168562 709392 168646 709628
rect 168882 709392 204326 709628
rect 204562 709392 204646 709628
rect 204882 709392 240326 709628
rect 240562 709392 240646 709628
rect 240882 709392 276326 709628
rect 276562 709392 276646 709628
rect 276882 709392 312326 709628
rect 312562 709392 312646 709628
rect 312882 709392 348326 709628
rect 348562 709392 348646 709628
rect 348882 709392 384326 709628
rect 384562 709392 384646 709628
rect 384882 709392 420326 709628
rect 420562 709392 420646 709628
rect 420882 709392 456326 709628
rect 456562 709392 456646 709628
rect 456882 709392 492326 709628
rect 492562 709392 492646 709628
rect 492882 709392 528326 709628
rect 528562 709392 528646 709628
rect 528882 709392 564326 709628
rect 564562 709392 564646 709628
rect 564882 709392 590452 709628
rect 590688 709392 590772 709628
rect 591008 709392 591040 709628
rect -7116 709360 591040 709392
rect -6156 708988 590080 709020
rect -6156 708752 -6124 708988
rect -5888 708752 -5804 708988
rect -5568 708752 19826 708988
rect 20062 708752 20146 708988
rect 20382 708752 55826 708988
rect 56062 708752 56146 708988
rect 56382 708752 91826 708988
rect 92062 708752 92146 708988
rect 92382 708752 127826 708988
rect 128062 708752 128146 708988
rect 128382 708752 163826 708988
rect 164062 708752 164146 708988
rect 164382 708752 199826 708988
rect 200062 708752 200146 708988
rect 200382 708752 235826 708988
rect 236062 708752 236146 708988
rect 236382 708752 271826 708988
rect 272062 708752 272146 708988
rect 272382 708752 307826 708988
rect 308062 708752 308146 708988
rect 308382 708752 343826 708988
rect 344062 708752 344146 708988
rect 344382 708752 379826 708988
rect 380062 708752 380146 708988
rect 380382 708752 415826 708988
rect 416062 708752 416146 708988
rect 416382 708752 451826 708988
rect 452062 708752 452146 708988
rect 452382 708752 487826 708988
rect 488062 708752 488146 708988
rect 488382 708752 523826 708988
rect 524062 708752 524146 708988
rect 524382 708752 559826 708988
rect 560062 708752 560146 708988
rect 560382 708752 589492 708988
rect 589728 708752 589812 708988
rect 590048 708752 590080 708988
rect -6156 708668 590080 708752
rect -6156 708432 -6124 708668
rect -5888 708432 -5804 708668
rect -5568 708432 19826 708668
rect 20062 708432 20146 708668
rect 20382 708432 55826 708668
rect 56062 708432 56146 708668
rect 56382 708432 91826 708668
rect 92062 708432 92146 708668
rect 92382 708432 127826 708668
rect 128062 708432 128146 708668
rect 128382 708432 163826 708668
rect 164062 708432 164146 708668
rect 164382 708432 199826 708668
rect 200062 708432 200146 708668
rect 200382 708432 235826 708668
rect 236062 708432 236146 708668
rect 236382 708432 271826 708668
rect 272062 708432 272146 708668
rect 272382 708432 307826 708668
rect 308062 708432 308146 708668
rect 308382 708432 343826 708668
rect 344062 708432 344146 708668
rect 344382 708432 379826 708668
rect 380062 708432 380146 708668
rect 380382 708432 415826 708668
rect 416062 708432 416146 708668
rect 416382 708432 451826 708668
rect 452062 708432 452146 708668
rect 452382 708432 487826 708668
rect 488062 708432 488146 708668
rect 488382 708432 523826 708668
rect 524062 708432 524146 708668
rect 524382 708432 559826 708668
rect 560062 708432 560146 708668
rect 560382 708432 589492 708668
rect 589728 708432 589812 708668
rect 590048 708432 590080 708668
rect -6156 708400 590080 708432
rect -5196 708028 589120 708060
rect -5196 707792 -5164 708028
rect -4928 707792 -4844 708028
rect -4608 707792 15326 708028
rect 15562 707792 15646 708028
rect 15882 707792 51326 708028
rect 51562 707792 51646 708028
rect 51882 707792 87326 708028
rect 87562 707792 87646 708028
rect 87882 707792 123326 708028
rect 123562 707792 123646 708028
rect 123882 707792 159326 708028
rect 159562 707792 159646 708028
rect 159882 707792 195326 708028
rect 195562 707792 195646 708028
rect 195882 707792 231326 708028
rect 231562 707792 231646 708028
rect 231882 707792 267326 708028
rect 267562 707792 267646 708028
rect 267882 707792 303326 708028
rect 303562 707792 303646 708028
rect 303882 707792 339326 708028
rect 339562 707792 339646 708028
rect 339882 707792 375326 708028
rect 375562 707792 375646 708028
rect 375882 707792 411326 708028
rect 411562 707792 411646 708028
rect 411882 707792 447326 708028
rect 447562 707792 447646 708028
rect 447882 707792 483326 708028
rect 483562 707792 483646 708028
rect 483882 707792 519326 708028
rect 519562 707792 519646 708028
rect 519882 707792 555326 708028
rect 555562 707792 555646 708028
rect 555882 707792 588532 708028
rect 588768 707792 588852 708028
rect 589088 707792 589120 708028
rect -5196 707708 589120 707792
rect -5196 707472 -5164 707708
rect -4928 707472 -4844 707708
rect -4608 707472 15326 707708
rect 15562 707472 15646 707708
rect 15882 707472 51326 707708
rect 51562 707472 51646 707708
rect 51882 707472 87326 707708
rect 87562 707472 87646 707708
rect 87882 707472 123326 707708
rect 123562 707472 123646 707708
rect 123882 707472 159326 707708
rect 159562 707472 159646 707708
rect 159882 707472 195326 707708
rect 195562 707472 195646 707708
rect 195882 707472 231326 707708
rect 231562 707472 231646 707708
rect 231882 707472 267326 707708
rect 267562 707472 267646 707708
rect 267882 707472 303326 707708
rect 303562 707472 303646 707708
rect 303882 707472 339326 707708
rect 339562 707472 339646 707708
rect 339882 707472 375326 707708
rect 375562 707472 375646 707708
rect 375882 707472 411326 707708
rect 411562 707472 411646 707708
rect 411882 707472 447326 707708
rect 447562 707472 447646 707708
rect 447882 707472 483326 707708
rect 483562 707472 483646 707708
rect 483882 707472 519326 707708
rect 519562 707472 519646 707708
rect 519882 707472 555326 707708
rect 555562 707472 555646 707708
rect 555882 707472 588532 707708
rect 588768 707472 588852 707708
rect 589088 707472 589120 707708
rect -5196 707440 589120 707472
rect -4236 707068 588160 707100
rect -4236 706832 -4204 707068
rect -3968 706832 -3884 707068
rect -3648 706832 10826 707068
rect 11062 706832 11146 707068
rect 11382 706832 46826 707068
rect 47062 706832 47146 707068
rect 47382 706832 82826 707068
rect 83062 706832 83146 707068
rect 83382 706832 118826 707068
rect 119062 706832 119146 707068
rect 119382 706832 154826 707068
rect 155062 706832 155146 707068
rect 155382 706832 190826 707068
rect 191062 706832 191146 707068
rect 191382 706832 226826 707068
rect 227062 706832 227146 707068
rect 227382 706832 262826 707068
rect 263062 706832 263146 707068
rect 263382 706832 298826 707068
rect 299062 706832 299146 707068
rect 299382 706832 334826 707068
rect 335062 706832 335146 707068
rect 335382 706832 370826 707068
rect 371062 706832 371146 707068
rect 371382 706832 406826 707068
rect 407062 706832 407146 707068
rect 407382 706832 442826 707068
rect 443062 706832 443146 707068
rect 443382 706832 478826 707068
rect 479062 706832 479146 707068
rect 479382 706832 514826 707068
rect 515062 706832 515146 707068
rect 515382 706832 550826 707068
rect 551062 706832 551146 707068
rect 551382 706832 587572 707068
rect 587808 706832 587892 707068
rect 588128 706832 588160 707068
rect -4236 706748 588160 706832
rect -4236 706512 -4204 706748
rect -3968 706512 -3884 706748
rect -3648 706512 10826 706748
rect 11062 706512 11146 706748
rect 11382 706512 46826 706748
rect 47062 706512 47146 706748
rect 47382 706512 82826 706748
rect 83062 706512 83146 706748
rect 83382 706512 118826 706748
rect 119062 706512 119146 706748
rect 119382 706512 154826 706748
rect 155062 706512 155146 706748
rect 155382 706512 190826 706748
rect 191062 706512 191146 706748
rect 191382 706512 226826 706748
rect 227062 706512 227146 706748
rect 227382 706512 262826 706748
rect 263062 706512 263146 706748
rect 263382 706512 298826 706748
rect 299062 706512 299146 706748
rect 299382 706512 334826 706748
rect 335062 706512 335146 706748
rect 335382 706512 370826 706748
rect 371062 706512 371146 706748
rect 371382 706512 406826 706748
rect 407062 706512 407146 706748
rect 407382 706512 442826 706748
rect 443062 706512 443146 706748
rect 443382 706512 478826 706748
rect 479062 706512 479146 706748
rect 479382 706512 514826 706748
rect 515062 706512 515146 706748
rect 515382 706512 550826 706748
rect 551062 706512 551146 706748
rect 551382 706512 587572 706748
rect 587808 706512 587892 706748
rect 588128 706512 588160 706748
rect -4236 706480 588160 706512
rect -3276 706108 587200 706140
rect -3276 705872 -3244 706108
rect -3008 705872 -2924 706108
rect -2688 705872 6326 706108
rect 6562 705872 6646 706108
rect 6882 705872 42326 706108
rect 42562 705872 42646 706108
rect 42882 705872 78326 706108
rect 78562 705872 78646 706108
rect 78882 705872 114326 706108
rect 114562 705872 114646 706108
rect 114882 705872 150326 706108
rect 150562 705872 150646 706108
rect 150882 705872 186326 706108
rect 186562 705872 186646 706108
rect 186882 705872 222326 706108
rect 222562 705872 222646 706108
rect 222882 705872 258326 706108
rect 258562 705872 258646 706108
rect 258882 705872 294326 706108
rect 294562 705872 294646 706108
rect 294882 705872 330326 706108
rect 330562 705872 330646 706108
rect 330882 705872 366326 706108
rect 366562 705872 366646 706108
rect 366882 705872 402326 706108
rect 402562 705872 402646 706108
rect 402882 705872 438326 706108
rect 438562 705872 438646 706108
rect 438882 705872 474326 706108
rect 474562 705872 474646 706108
rect 474882 705872 510326 706108
rect 510562 705872 510646 706108
rect 510882 705872 546326 706108
rect 546562 705872 546646 706108
rect 546882 705872 582326 706108
rect 582562 705872 582646 706108
rect 582882 705872 586612 706108
rect 586848 705872 586932 706108
rect 587168 705872 587200 706108
rect -3276 705788 587200 705872
rect -3276 705552 -3244 705788
rect -3008 705552 -2924 705788
rect -2688 705552 6326 705788
rect 6562 705552 6646 705788
rect 6882 705552 42326 705788
rect 42562 705552 42646 705788
rect 42882 705552 78326 705788
rect 78562 705552 78646 705788
rect 78882 705552 114326 705788
rect 114562 705552 114646 705788
rect 114882 705552 150326 705788
rect 150562 705552 150646 705788
rect 150882 705552 186326 705788
rect 186562 705552 186646 705788
rect 186882 705552 222326 705788
rect 222562 705552 222646 705788
rect 222882 705552 258326 705788
rect 258562 705552 258646 705788
rect 258882 705552 294326 705788
rect 294562 705552 294646 705788
rect 294882 705552 330326 705788
rect 330562 705552 330646 705788
rect 330882 705552 366326 705788
rect 366562 705552 366646 705788
rect 366882 705552 402326 705788
rect 402562 705552 402646 705788
rect 402882 705552 438326 705788
rect 438562 705552 438646 705788
rect 438882 705552 474326 705788
rect 474562 705552 474646 705788
rect 474882 705552 510326 705788
rect 510562 705552 510646 705788
rect 510882 705552 546326 705788
rect 546562 705552 546646 705788
rect 546882 705552 582326 705788
rect 582562 705552 582646 705788
rect 582882 705552 586612 705788
rect 586848 705552 586932 705788
rect 587168 705552 587200 705788
rect -3276 705520 587200 705552
rect -2316 705148 586240 705180
rect -2316 704912 -2284 705148
rect -2048 704912 -1964 705148
rect -1728 704912 1826 705148
rect 2062 704912 2146 705148
rect 2382 704912 37826 705148
rect 38062 704912 38146 705148
rect 38382 704912 73826 705148
rect 74062 704912 74146 705148
rect 74382 704912 109826 705148
rect 110062 704912 110146 705148
rect 110382 704912 145826 705148
rect 146062 704912 146146 705148
rect 146382 704912 181826 705148
rect 182062 704912 182146 705148
rect 182382 704912 217826 705148
rect 218062 704912 218146 705148
rect 218382 704912 253826 705148
rect 254062 704912 254146 705148
rect 254382 704912 289826 705148
rect 290062 704912 290146 705148
rect 290382 704912 325826 705148
rect 326062 704912 326146 705148
rect 326382 704912 361826 705148
rect 362062 704912 362146 705148
rect 362382 704912 397826 705148
rect 398062 704912 398146 705148
rect 398382 704912 433826 705148
rect 434062 704912 434146 705148
rect 434382 704912 469826 705148
rect 470062 704912 470146 705148
rect 470382 704912 505826 705148
rect 506062 704912 506146 705148
rect 506382 704912 541826 705148
rect 542062 704912 542146 705148
rect 542382 704912 577826 705148
rect 578062 704912 578146 705148
rect 578382 704912 585652 705148
rect 585888 704912 585972 705148
rect 586208 704912 586240 705148
rect -2316 704828 586240 704912
rect -2316 704592 -2284 704828
rect -2048 704592 -1964 704828
rect -1728 704592 1826 704828
rect 2062 704592 2146 704828
rect 2382 704592 37826 704828
rect 38062 704592 38146 704828
rect 38382 704592 73826 704828
rect 74062 704592 74146 704828
rect 74382 704592 109826 704828
rect 110062 704592 110146 704828
rect 110382 704592 145826 704828
rect 146062 704592 146146 704828
rect 146382 704592 181826 704828
rect 182062 704592 182146 704828
rect 182382 704592 217826 704828
rect 218062 704592 218146 704828
rect 218382 704592 253826 704828
rect 254062 704592 254146 704828
rect 254382 704592 289826 704828
rect 290062 704592 290146 704828
rect 290382 704592 325826 704828
rect 326062 704592 326146 704828
rect 326382 704592 361826 704828
rect 362062 704592 362146 704828
rect 362382 704592 397826 704828
rect 398062 704592 398146 704828
rect 398382 704592 433826 704828
rect 434062 704592 434146 704828
rect 434382 704592 469826 704828
rect 470062 704592 470146 704828
rect 470382 704592 505826 704828
rect 506062 704592 506146 704828
rect 506382 704592 541826 704828
rect 542062 704592 542146 704828
rect 542382 704592 577826 704828
rect 578062 704592 578146 704828
rect 578382 704592 585652 704828
rect 585888 704592 585972 704828
rect 586208 704592 586240 704828
rect -2316 704560 586240 704592
rect -9036 700954 592960 700986
rect -9036 700718 -5164 700954
rect -4928 700718 -4844 700954
rect -4608 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588532 700954
rect 588768 700718 588852 700954
rect 589088 700718 592960 700954
rect -9036 700634 592960 700718
rect -9036 700398 -5164 700634
rect -4928 700398 -4844 700634
rect -4608 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588532 700634
rect 588768 700398 588852 700634
rect 589088 700398 592960 700634
rect -9036 700366 592960 700398
rect -9036 696454 592960 696486
rect -9036 696218 -4204 696454
rect -3968 696218 -3884 696454
rect -3648 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587572 696454
rect 587808 696218 587892 696454
rect 588128 696218 592960 696454
rect -9036 696134 592960 696218
rect -9036 695898 -4204 696134
rect -3968 695898 -3884 696134
rect -3648 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587572 696134
rect 587808 695898 587892 696134
rect 588128 695898 592960 696134
rect -9036 695866 592960 695898
rect -9036 691954 592960 691986
rect -9036 691718 -3244 691954
rect -3008 691718 -2924 691954
rect -2688 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586612 691954
rect 586848 691718 586932 691954
rect 587168 691718 592960 691954
rect -9036 691634 592960 691718
rect -9036 691398 -3244 691634
rect -3008 691398 -2924 691634
rect -2688 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586612 691634
rect 586848 691398 586932 691634
rect 587168 691398 592960 691634
rect -9036 691366 592960 691398
rect -9036 687454 592960 687486
rect -9036 687218 -2284 687454
rect -2048 687218 -1964 687454
rect -1728 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585652 687454
rect 585888 687218 585972 687454
rect 586208 687218 592960 687454
rect -9036 687134 592960 687218
rect -9036 686898 -2284 687134
rect -2048 686898 -1964 687134
rect -1728 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585652 687134
rect 585888 686898 585972 687134
rect 586208 686898 592960 687134
rect -9036 686866 592960 686898
rect -9036 682954 592960 682986
rect -9036 682718 -9004 682954
rect -8768 682718 -8684 682954
rect -8448 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592372 682954
rect 592608 682718 592692 682954
rect 592928 682718 592960 682954
rect -9036 682634 592960 682718
rect -9036 682398 -9004 682634
rect -8768 682398 -8684 682634
rect -8448 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592372 682634
rect 592608 682398 592692 682634
rect 592928 682398 592960 682634
rect -9036 682366 592960 682398
rect -9036 678454 592960 678486
rect -9036 678218 -8044 678454
rect -7808 678218 -7724 678454
rect -7488 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591412 678454
rect 591648 678218 591732 678454
rect 591968 678218 592960 678454
rect -9036 678134 592960 678218
rect -9036 677898 -8044 678134
rect -7808 677898 -7724 678134
rect -7488 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591412 678134
rect 591648 677898 591732 678134
rect 591968 677898 592960 678134
rect -9036 677866 592960 677898
rect -9036 673954 592960 673986
rect -9036 673718 -7084 673954
rect -6848 673718 -6764 673954
rect -6528 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590452 673954
rect 590688 673718 590772 673954
rect 591008 673718 592960 673954
rect -9036 673634 592960 673718
rect -9036 673398 -7084 673634
rect -6848 673398 -6764 673634
rect -6528 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590452 673634
rect 590688 673398 590772 673634
rect 591008 673398 592960 673634
rect -9036 673366 592960 673398
rect -9036 669454 592960 669486
rect -9036 669218 -6124 669454
rect -5888 669218 -5804 669454
rect -5568 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589492 669454
rect 589728 669218 589812 669454
rect 590048 669218 592960 669454
rect -9036 669134 592960 669218
rect -9036 668898 -6124 669134
rect -5888 668898 -5804 669134
rect -5568 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589492 669134
rect 589728 668898 589812 669134
rect 590048 668898 592960 669134
rect -9036 668866 592960 668898
rect -9036 664954 592960 664986
rect -9036 664718 -5164 664954
rect -4928 664718 -4844 664954
rect -4608 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588532 664954
rect 588768 664718 588852 664954
rect 589088 664718 592960 664954
rect -9036 664634 592960 664718
rect -9036 664398 -5164 664634
rect -4928 664398 -4844 664634
rect -4608 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588532 664634
rect 588768 664398 588852 664634
rect 589088 664398 592960 664634
rect -9036 664366 592960 664398
rect -9036 660454 592960 660486
rect -9036 660218 -4204 660454
rect -3968 660218 -3884 660454
rect -3648 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587572 660454
rect 587808 660218 587892 660454
rect 588128 660218 592960 660454
rect -9036 660134 592960 660218
rect -9036 659898 -4204 660134
rect -3968 659898 -3884 660134
rect -3648 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587572 660134
rect 587808 659898 587892 660134
rect 588128 659898 592960 660134
rect -9036 659866 592960 659898
rect -9036 655954 592960 655986
rect -9036 655718 -3244 655954
rect -3008 655718 -2924 655954
rect -2688 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586612 655954
rect 586848 655718 586932 655954
rect 587168 655718 592960 655954
rect -9036 655634 592960 655718
rect -9036 655398 -3244 655634
rect -3008 655398 -2924 655634
rect -2688 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586612 655634
rect 586848 655398 586932 655634
rect 587168 655398 592960 655634
rect -9036 655366 592960 655398
rect -9036 651454 592960 651486
rect -9036 651218 -2284 651454
rect -2048 651218 -1964 651454
rect -1728 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585652 651454
rect 585888 651218 585972 651454
rect 586208 651218 592960 651454
rect -9036 651134 592960 651218
rect -9036 650898 -2284 651134
rect -2048 650898 -1964 651134
rect -1728 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585652 651134
rect 585888 650898 585972 651134
rect 586208 650898 592960 651134
rect -9036 650866 592960 650898
rect -9036 646954 592960 646986
rect -9036 646718 -9004 646954
rect -8768 646718 -8684 646954
rect -8448 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592372 646954
rect 592608 646718 592692 646954
rect 592928 646718 592960 646954
rect -9036 646634 592960 646718
rect -9036 646398 -9004 646634
rect -8768 646398 -8684 646634
rect -8448 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592372 646634
rect 592608 646398 592692 646634
rect 592928 646398 592960 646634
rect -9036 646366 592960 646398
rect -9036 642454 592960 642486
rect -9036 642218 -8044 642454
rect -7808 642218 -7724 642454
rect -7488 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591412 642454
rect 591648 642218 591732 642454
rect 591968 642218 592960 642454
rect -9036 642134 592960 642218
rect -9036 641898 -8044 642134
rect -7808 641898 -7724 642134
rect -7488 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591412 642134
rect 591648 641898 591732 642134
rect 591968 641898 592960 642134
rect -9036 641866 592960 641898
rect -9036 637954 592960 637986
rect -9036 637718 -7084 637954
rect -6848 637718 -6764 637954
rect -6528 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590452 637954
rect 590688 637718 590772 637954
rect 591008 637718 592960 637954
rect -9036 637634 592960 637718
rect -9036 637398 -7084 637634
rect -6848 637398 -6764 637634
rect -6528 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590452 637634
rect 590688 637398 590772 637634
rect 591008 637398 592960 637634
rect -9036 637366 592960 637398
rect -9036 633454 592960 633486
rect -9036 633218 -6124 633454
rect -5888 633218 -5804 633454
rect -5568 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589492 633454
rect 589728 633218 589812 633454
rect 590048 633218 592960 633454
rect -9036 633134 592960 633218
rect -9036 632898 -6124 633134
rect -5888 632898 -5804 633134
rect -5568 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589492 633134
rect 589728 632898 589812 633134
rect 590048 632898 592960 633134
rect -9036 632866 592960 632898
rect -9036 628954 592960 628986
rect -9036 628718 -5164 628954
rect -4928 628718 -4844 628954
rect -4608 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588532 628954
rect 588768 628718 588852 628954
rect 589088 628718 592960 628954
rect -9036 628634 592960 628718
rect -9036 628398 -5164 628634
rect -4928 628398 -4844 628634
rect -4608 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588532 628634
rect 588768 628398 588852 628634
rect 589088 628398 592960 628634
rect -9036 628366 592960 628398
rect -9036 624454 592960 624486
rect -9036 624218 -4204 624454
rect -3968 624218 -3884 624454
rect -3648 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587572 624454
rect 587808 624218 587892 624454
rect 588128 624218 592960 624454
rect -9036 624134 592960 624218
rect -9036 623898 -4204 624134
rect -3968 623898 -3884 624134
rect -3648 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587572 624134
rect 587808 623898 587892 624134
rect 588128 623898 592960 624134
rect -9036 623866 592960 623898
rect -9036 619954 592960 619986
rect -9036 619718 -3244 619954
rect -3008 619718 -2924 619954
rect -2688 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586612 619954
rect 586848 619718 586932 619954
rect 587168 619718 592960 619954
rect -9036 619634 592960 619718
rect -9036 619398 -3244 619634
rect -3008 619398 -2924 619634
rect -2688 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586612 619634
rect 586848 619398 586932 619634
rect 587168 619398 592960 619634
rect -9036 619366 592960 619398
rect -9036 615454 592960 615486
rect -9036 615218 -2284 615454
rect -2048 615218 -1964 615454
rect -1728 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585652 615454
rect 585888 615218 585972 615454
rect 586208 615218 592960 615454
rect -9036 615134 592960 615218
rect -9036 614898 -2284 615134
rect -2048 614898 -1964 615134
rect -1728 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585652 615134
rect 585888 614898 585972 615134
rect 586208 614898 592960 615134
rect -9036 614866 592960 614898
rect -9036 610954 592960 610986
rect -9036 610718 -9004 610954
rect -8768 610718 -8684 610954
rect -8448 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592372 610954
rect 592608 610718 592692 610954
rect 592928 610718 592960 610954
rect -9036 610634 592960 610718
rect -9036 610398 -9004 610634
rect -8768 610398 -8684 610634
rect -8448 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592372 610634
rect 592608 610398 592692 610634
rect 592928 610398 592960 610634
rect -9036 610366 592960 610398
rect -9036 606454 592960 606486
rect -9036 606218 -8044 606454
rect -7808 606218 -7724 606454
rect -7488 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591412 606454
rect 591648 606218 591732 606454
rect 591968 606218 592960 606454
rect -9036 606134 592960 606218
rect -9036 605898 -8044 606134
rect -7808 605898 -7724 606134
rect -7488 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591412 606134
rect 591648 605898 591732 606134
rect 591968 605898 592960 606134
rect -9036 605866 592960 605898
rect -9036 601954 592960 601986
rect -9036 601718 -7084 601954
rect -6848 601718 -6764 601954
rect -6528 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590452 601954
rect 590688 601718 590772 601954
rect 591008 601718 592960 601954
rect -9036 601634 592960 601718
rect -9036 601398 -7084 601634
rect -6848 601398 -6764 601634
rect -6528 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590452 601634
rect 590688 601398 590772 601634
rect 591008 601398 592960 601634
rect -9036 601366 592960 601398
rect -9036 597454 592960 597486
rect -9036 597218 -6124 597454
rect -5888 597218 -5804 597454
rect -5568 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589492 597454
rect 589728 597218 589812 597454
rect 590048 597218 592960 597454
rect -9036 597134 592960 597218
rect -9036 596898 -6124 597134
rect -5888 596898 -5804 597134
rect -5568 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589492 597134
rect 589728 596898 589812 597134
rect 590048 596898 592960 597134
rect -9036 596866 592960 596898
rect -9036 592954 592960 592986
rect -9036 592718 -5164 592954
rect -4928 592718 -4844 592954
rect -4608 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588532 592954
rect 588768 592718 588852 592954
rect 589088 592718 592960 592954
rect -9036 592634 592960 592718
rect -9036 592398 -5164 592634
rect -4928 592398 -4844 592634
rect -4608 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588532 592634
rect 588768 592398 588852 592634
rect 589088 592398 592960 592634
rect -9036 592366 592960 592398
rect -9036 588454 592960 588486
rect -9036 588218 -4204 588454
rect -3968 588218 -3884 588454
rect -3648 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587572 588454
rect 587808 588218 587892 588454
rect 588128 588218 592960 588454
rect -9036 588134 592960 588218
rect -9036 587898 -4204 588134
rect -3968 587898 -3884 588134
rect -3648 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587572 588134
rect 587808 587898 587892 588134
rect 588128 587898 592960 588134
rect -9036 587866 592960 587898
rect -9036 583954 592960 583986
rect -9036 583718 -3244 583954
rect -3008 583718 -2924 583954
rect -2688 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586612 583954
rect 586848 583718 586932 583954
rect 587168 583718 592960 583954
rect -9036 583634 592960 583718
rect -9036 583398 -3244 583634
rect -3008 583398 -2924 583634
rect -2688 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586612 583634
rect 586848 583398 586932 583634
rect 587168 583398 592960 583634
rect -9036 583366 592960 583398
rect -9036 579454 592960 579486
rect -9036 579218 -2284 579454
rect -2048 579218 -1964 579454
rect -1728 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585652 579454
rect 585888 579218 585972 579454
rect 586208 579218 592960 579454
rect -9036 579134 592960 579218
rect -9036 578898 -2284 579134
rect -2048 578898 -1964 579134
rect -1728 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585652 579134
rect 585888 578898 585972 579134
rect 586208 578898 592960 579134
rect -9036 578866 592960 578898
rect -9036 574954 592960 574986
rect -9036 574718 -9004 574954
rect -8768 574718 -8684 574954
rect -8448 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592372 574954
rect 592608 574718 592692 574954
rect 592928 574718 592960 574954
rect -9036 574634 592960 574718
rect -9036 574398 -9004 574634
rect -8768 574398 -8684 574634
rect -8448 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592372 574634
rect 592608 574398 592692 574634
rect 592928 574398 592960 574634
rect -9036 574366 592960 574398
rect -9036 570454 592960 570486
rect -9036 570218 -8044 570454
rect -7808 570218 -7724 570454
rect -7488 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591412 570454
rect 591648 570218 591732 570454
rect 591968 570218 592960 570454
rect -9036 570134 592960 570218
rect -9036 569898 -8044 570134
rect -7808 569898 -7724 570134
rect -7488 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591412 570134
rect 591648 569898 591732 570134
rect 591968 569898 592960 570134
rect -9036 569866 592960 569898
rect -9036 565954 592960 565986
rect -9036 565718 -7084 565954
rect -6848 565718 -6764 565954
rect -6528 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590452 565954
rect 590688 565718 590772 565954
rect 591008 565718 592960 565954
rect -9036 565634 592960 565718
rect -9036 565398 -7084 565634
rect -6848 565398 -6764 565634
rect -6528 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590452 565634
rect 590688 565398 590772 565634
rect 591008 565398 592960 565634
rect -9036 565366 592960 565398
rect -9036 561454 592960 561486
rect -9036 561218 -6124 561454
rect -5888 561218 -5804 561454
rect -5568 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589492 561454
rect 589728 561218 589812 561454
rect 590048 561218 592960 561454
rect -9036 561134 592960 561218
rect -9036 560898 -6124 561134
rect -5888 560898 -5804 561134
rect -5568 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589492 561134
rect 589728 560898 589812 561134
rect 590048 560898 592960 561134
rect -9036 560866 592960 560898
rect -9036 556954 592960 556986
rect -9036 556718 -5164 556954
rect -4928 556718 -4844 556954
rect -4608 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588532 556954
rect 588768 556718 588852 556954
rect 589088 556718 592960 556954
rect -9036 556634 592960 556718
rect -9036 556398 -5164 556634
rect -4928 556398 -4844 556634
rect -4608 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588532 556634
rect 588768 556398 588852 556634
rect 589088 556398 592960 556634
rect -9036 556366 592960 556398
rect -9036 552454 592960 552486
rect -9036 552218 -4204 552454
rect -3968 552218 -3884 552454
rect -3648 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587572 552454
rect 587808 552218 587892 552454
rect 588128 552218 592960 552454
rect -9036 552134 592960 552218
rect -9036 551898 -4204 552134
rect -3968 551898 -3884 552134
rect -3648 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587572 552134
rect 587808 551898 587892 552134
rect 588128 551898 592960 552134
rect -9036 551866 592960 551898
rect -9036 547954 592960 547986
rect -9036 547718 -3244 547954
rect -3008 547718 -2924 547954
rect -2688 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586612 547954
rect 586848 547718 586932 547954
rect 587168 547718 592960 547954
rect -9036 547634 592960 547718
rect -9036 547398 -3244 547634
rect -3008 547398 -2924 547634
rect -2688 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586612 547634
rect 586848 547398 586932 547634
rect 587168 547398 592960 547634
rect -9036 547366 592960 547398
rect -9036 543454 592960 543486
rect -9036 543218 -2284 543454
rect -2048 543218 -1964 543454
rect -1728 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585652 543454
rect 585888 543218 585972 543454
rect 586208 543218 592960 543454
rect -9036 543134 592960 543218
rect -9036 542898 -2284 543134
rect -2048 542898 -1964 543134
rect -1728 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585652 543134
rect 585888 542898 585972 543134
rect 586208 542898 592960 543134
rect -9036 542866 592960 542898
rect -9036 538954 592960 538986
rect -9036 538718 -9004 538954
rect -8768 538718 -8684 538954
rect -8448 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592372 538954
rect 592608 538718 592692 538954
rect 592928 538718 592960 538954
rect -9036 538634 592960 538718
rect -9036 538398 -9004 538634
rect -8768 538398 -8684 538634
rect -8448 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592372 538634
rect 592608 538398 592692 538634
rect 592928 538398 592960 538634
rect -9036 538366 592960 538398
rect -9036 534454 592960 534486
rect -9036 534218 -8044 534454
rect -7808 534218 -7724 534454
rect -7488 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591412 534454
rect 591648 534218 591732 534454
rect 591968 534218 592960 534454
rect -9036 534134 592960 534218
rect -9036 533898 -8044 534134
rect -7808 533898 -7724 534134
rect -7488 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591412 534134
rect 591648 533898 591732 534134
rect 591968 533898 592960 534134
rect -9036 533866 592960 533898
rect -9036 529954 592960 529986
rect -9036 529718 -7084 529954
rect -6848 529718 -6764 529954
rect -6528 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590452 529954
rect 590688 529718 590772 529954
rect 591008 529718 592960 529954
rect -9036 529634 592960 529718
rect -9036 529398 -7084 529634
rect -6848 529398 -6764 529634
rect -6528 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590452 529634
rect 590688 529398 590772 529634
rect 591008 529398 592960 529634
rect -9036 529366 592960 529398
rect -9036 525454 592960 525486
rect -9036 525218 -6124 525454
rect -5888 525218 -5804 525454
rect -5568 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589492 525454
rect 589728 525218 589812 525454
rect 590048 525218 592960 525454
rect -9036 525134 592960 525218
rect -9036 524898 -6124 525134
rect -5888 524898 -5804 525134
rect -5568 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589492 525134
rect 589728 524898 589812 525134
rect 590048 524898 592960 525134
rect -9036 524866 592960 524898
rect -9036 520954 592960 520986
rect -9036 520718 -5164 520954
rect -4928 520718 -4844 520954
rect -4608 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588532 520954
rect 588768 520718 588852 520954
rect 589088 520718 592960 520954
rect -9036 520634 592960 520718
rect -9036 520398 -5164 520634
rect -4928 520398 -4844 520634
rect -4608 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588532 520634
rect 588768 520398 588852 520634
rect 589088 520398 592960 520634
rect -9036 520366 592960 520398
rect -9036 516454 592960 516486
rect -9036 516218 -4204 516454
rect -3968 516218 -3884 516454
rect -3648 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587572 516454
rect 587808 516218 587892 516454
rect 588128 516218 592960 516454
rect -9036 516134 592960 516218
rect -9036 515898 -4204 516134
rect -3968 515898 -3884 516134
rect -3648 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587572 516134
rect 587808 515898 587892 516134
rect 588128 515898 592960 516134
rect -9036 515866 592960 515898
rect -9036 511954 592960 511986
rect -9036 511718 -3244 511954
rect -3008 511718 -2924 511954
rect -2688 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586612 511954
rect 586848 511718 586932 511954
rect 587168 511718 592960 511954
rect -9036 511634 592960 511718
rect -9036 511398 -3244 511634
rect -3008 511398 -2924 511634
rect -2688 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586612 511634
rect 586848 511398 586932 511634
rect 587168 511398 592960 511634
rect -9036 511366 592960 511398
rect -9036 507454 592960 507486
rect -9036 507218 -2284 507454
rect -2048 507218 -1964 507454
rect -1728 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585652 507454
rect 585888 507218 585972 507454
rect 586208 507218 592960 507454
rect -9036 507134 592960 507218
rect -9036 506898 -2284 507134
rect -2048 506898 -1964 507134
rect -1728 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585652 507134
rect 585888 506898 585972 507134
rect 586208 506898 592960 507134
rect -9036 506866 592960 506898
rect -9036 502954 592960 502986
rect -9036 502718 -9004 502954
rect -8768 502718 -8684 502954
rect -8448 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592372 502954
rect 592608 502718 592692 502954
rect 592928 502718 592960 502954
rect -9036 502634 592960 502718
rect -9036 502398 -9004 502634
rect -8768 502398 -8684 502634
rect -8448 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592372 502634
rect 592608 502398 592692 502634
rect 592928 502398 592960 502634
rect -9036 502366 592960 502398
rect -9036 498454 592960 498486
rect -9036 498218 -8044 498454
rect -7808 498218 -7724 498454
rect -7488 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591412 498454
rect 591648 498218 591732 498454
rect 591968 498218 592960 498454
rect -9036 498134 592960 498218
rect -9036 497898 -8044 498134
rect -7808 497898 -7724 498134
rect -7488 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591412 498134
rect 591648 497898 591732 498134
rect 591968 497898 592960 498134
rect -9036 497866 592960 497898
rect -9036 493954 592960 493986
rect -9036 493718 -7084 493954
rect -6848 493718 -6764 493954
rect -6528 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590452 493954
rect 590688 493718 590772 493954
rect 591008 493718 592960 493954
rect -9036 493634 592960 493718
rect -9036 493398 -7084 493634
rect -6848 493398 -6764 493634
rect -6528 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590452 493634
rect 590688 493398 590772 493634
rect 591008 493398 592960 493634
rect -9036 493366 592960 493398
rect -9036 489454 592960 489486
rect -9036 489218 -6124 489454
rect -5888 489218 -5804 489454
rect -5568 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589492 489454
rect 589728 489218 589812 489454
rect 590048 489218 592960 489454
rect -9036 489134 592960 489218
rect -9036 488898 -6124 489134
rect -5888 488898 -5804 489134
rect -5568 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589492 489134
rect 589728 488898 589812 489134
rect 590048 488898 592960 489134
rect -9036 488866 592960 488898
rect -9036 484954 592960 484986
rect -9036 484718 -5164 484954
rect -4928 484718 -4844 484954
rect -4608 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588532 484954
rect 588768 484718 588852 484954
rect 589088 484718 592960 484954
rect -9036 484634 592960 484718
rect -9036 484398 -5164 484634
rect -4928 484398 -4844 484634
rect -4608 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588532 484634
rect 588768 484398 588852 484634
rect 589088 484398 592960 484634
rect -9036 484366 592960 484398
rect -9036 480454 592960 480486
rect -9036 480218 -4204 480454
rect -3968 480218 -3884 480454
rect -3648 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587572 480454
rect 587808 480218 587892 480454
rect 588128 480218 592960 480454
rect -9036 480134 592960 480218
rect -9036 479898 -4204 480134
rect -3968 479898 -3884 480134
rect -3648 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587572 480134
rect 587808 479898 587892 480134
rect 588128 479898 592960 480134
rect -9036 479866 592960 479898
rect -9036 475954 592960 475986
rect -9036 475718 -3244 475954
rect -3008 475718 -2924 475954
rect -2688 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586612 475954
rect 586848 475718 586932 475954
rect 587168 475718 592960 475954
rect -9036 475634 592960 475718
rect -9036 475398 -3244 475634
rect -3008 475398 -2924 475634
rect -2688 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586612 475634
rect 586848 475398 586932 475634
rect 587168 475398 592960 475634
rect -9036 475366 592960 475398
rect -9036 471454 592960 471486
rect -9036 471218 -2284 471454
rect -2048 471218 -1964 471454
rect -1728 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585652 471454
rect 585888 471218 585972 471454
rect 586208 471218 592960 471454
rect -9036 471134 592960 471218
rect -9036 470898 -2284 471134
rect -2048 470898 -1964 471134
rect -1728 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585652 471134
rect 585888 470898 585972 471134
rect 586208 470898 592960 471134
rect -9036 470866 592960 470898
rect -9036 466954 592960 466986
rect -9036 466718 -9004 466954
rect -8768 466718 -8684 466954
rect -8448 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592372 466954
rect 592608 466718 592692 466954
rect 592928 466718 592960 466954
rect -9036 466634 592960 466718
rect -9036 466398 -9004 466634
rect -8768 466398 -8684 466634
rect -8448 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592372 466634
rect 592608 466398 592692 466634
rect 592928 466398 592960 466634
rect -9036 466366 592960 466398
rect -9036 462454 592960 462486
rect -9036 462218 -8044 462454
rect -7808 462218 -7724 462454
rect -7488 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591412 462454
rect 591648 462218 591732 462454
rect 591968 462218 592960 462454
rect -9036 462134 592960 462218
rect -9036 461898 -8044 462134
rect -7808 461898 -7724 462134
rect -7488 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591412 462134
rect 591648 461898 591732 462134
rect 591968 461898 592960 462134
rect -9036 461866 592960 461898
rect -9036 457954 592960 457986
rect -9036 457718 -7084 457954
rect -6848 457718 -6764 457954
rect -6528 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590452 457954
rect 590688 457718 590772 457954
rect 591008 457718 592960 457954
rect -9036 457634 592960 457718
rect -9036 457398 -7084 457634
rect -6848 457398 -6764 457634
rect -6528 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590452 457634
rect 590688 457398 590772 457634
rect 591008 457398 592960 457634
rect -9036 457366 592960 457398
rect -9036 453454 592960 453486
rect -9036 453218 -6124 453454
rect -5888 453218 -5804 453454
rect -5568 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589492 453454
rect 589728 453218 589812 453454
rect 590048 453218 592960 453454
rect -9036 453134 592960 453218
rect -9036 452898 -6124 453134
rect -5888 452898 -5804 453134
rect -5568 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589492 453134
rect 589728 452898 589812 453134
rect 590048 452898 592960 453134
rect -9036 452866 592960 452898
rect -9036 448954 592960 448986
rect -9036 448718 -5164 448954
rect -4928 448718 -4844 448954
rect -4608 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588532 448954
rect 588768 448718 588852 448954
rect 589088 448718 592960 448954
rect -9036 448634 592960 448718
rect -9036 448398 -5164 448634
rect -4928 448398 -4844 448634
rect -4608 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588532 448634
rect 588768 448398 588852 448634
rect 589088 448398 592960 448634
rect -9036 448366 592960 448398
rect -9036 444454 592960 444486
rect -9036 444218 -4204 444454
rect -3968 444218 -3884 444454
rect -3648 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587572 444454
rect 587808 444218 587892 444454
rect 588128 444218 592960 444454
rect -9036 444134 592960 444218
rect -9036 443898 -4204 444134
rect -3968 443898 -3884 444134
rect -3648 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587572 444134
rect 587808 443898 587892 444134
rect 588128 443898 592960 444134
rect -9036 443866 592960 443898
rect -9036 439954 592960 439986
rect -9036 439718 -3244 439954
rect -3008 439718 -2924 439954
rect -2688 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586612 439954
rect 586848 439718 586932 439954
rect 587168 439718 592960 439954
rect -9036 439634 592960 439718
rect -9036 439398 -3244 439634
rect -3008 439398 -2924 439634
rect -2688 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586612 439634
rect 586848 439398 586932 439634
rect 587168 439398 592960 439634
rect -9036 439366 592960 439398
rect -9036 435454 592960 435486
rect -9036 435218 -2284 435454
rect -2048 435218 -1964 435454
rect -1728 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585652 435454
rect 585888 435218 585972 435454
rect 586208 435218 592960 435454
rect -9036 435134 592960 435218
rect -9036 434898 -2284 435134
rect -2048 434898 -1964 435134
rect -1728 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585652 435134
rect 585888 434898 585972 435134
rect 586208 434898 592960 435134
rect -9036 434866 592960 434898
rect -9036 430954 592960 430986
rect -9036 430718 -9004 430954
rect -8768 430718 -8684 430954
rect -8448 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592372 430954
rect 592608 430718 592692 430954
rect 592928 430718 592960 430954
rect -9036 430634 592960 430718
rect -9036 430398 -9004 430634
rect -8768 430398 -8684 430634
rect -8448 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592372 430634
rect 592608 430398 592692 430634
rect 592928 430398 592960 430634
rect -9036 430366 592960 430398
rect -9036 426454 592960 426486
rect -9036 426218 -8044 426454
rect -7808 426218 -7724 426454
rect -7488 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591412 426454
rect 591648 426218 591732 426454
rect 591968 426218 592960 426454
rect -9036 426134 592960 426218
rect -9036 425898 -8044 426134
rect -7808 425898 -7724 426134
rect -7488 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591412 426134
rect 591648 425898 591732 426134
rect 591968 425898 592960 426134
rect -9036 425866 592960 425898
rect -9036 421954 592960 421986
rect -9036 421718 -7084 421954
rect -6848 421718 -6764 421954
rect -6528 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590452 421954
rect 590688 421718 590772 421954
rect 591008 421718 592960 421954
rect -9036 421634 592960 421718
rect -9036 421398 -7084 421634
rect -6848 421398 -6764 421634
rect -6528 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590452 421634
rect 590688 421398 590772 421634
rect 591008 421398 592960 421634
rect -9036 421366 592960 421398
rect -9036 417454 592960 417486
rect -9036 417218 -6124 417454
rect -5888 417218 -5804 417454
rect -5568 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589492 417454
rect 589728 417218 589812 417454
rect 590048 417218 592960 417454
rect -9036 417134 592960 417218
rect -9036 416898 -6124 417134
rect -5888 416898 -5804 417134
rect -5568 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589492 417134
rect 589728 416898 589812 417134
rect 590048 416898 592960 417134
rect -9036 416866 592960 416898
rect -9036 412954 592960 412986
rect -9036 412718 -5164 412954
rect -4928 412718 -4844 412954
rect -4608 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588532 412954
rect 588768 412718 588852 412954
rect 589088 412718 592960 412954
rect -9036 412634 592960 412718
rect -9036 412398 -5164 412634
rect -4928 412398 -4844 412634
rect -4608 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588532 412634
rect 588768 412398 588852 412634
rect 589088 412398 592960 412634
rect -9036 412366 592960 412398
rect -9036 408454 592960 408486
rect -9036 408218 -4204 408454
rect -3968 408218 -3884 408454
rect -3648 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587572 408454
rect 587808 408218 587892 408454
rect 588128 408218 592960 408454
rect -9036 408134 592960 408218
rect -9036 407898 -4204 408134
rect -3968 407898 -3884 408134
rect -3648 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587572 408134
rect 587808 407898 587892 408134
rect 588128 407898 592960 408134
rect -9036 407866 592960 407898
rect -9036 403954 592960 403986
rect -9036 403718 -3244 403954
rect -3008 403718 -2924 403954
rect -2688 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586612 403954
rect 586848 403718 586932 403954
rect 587168 403718 592960 403954
rect -9036 403634 592960 403718
rect -9036 403398 -3244 403634
rect -3008 403398 -2924 403634
rect -2688 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586612 403634
rect 586848 403398 586932 403634
rect 587168 403398 592960 403634
rect -9036 403366 592960 403398
rect -9036 399454 592960 399486
rect -9036 399218 -2284 399454
rect -2048 399218 -1964 399454
rect -1728 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585652 399454
rect 585888 399218 585972 399454
rect 586208 399218 592960 399454
rect -9036 399134 592960 399218
rect -9036 398898 -2284 399134
rect -2048 398898 -1964 399134
rect -1728 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585652 399134
rect 585888 398898 585972 399134
rect 586208 398898 592960 399134
rect -9036 398866 592960 398898
rect -9036 394954 592960 394986
rect -9036 394718 -9004 394954
rect -8768 394718 -8684 394954
rect -8448 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592372 394954
rect 592608 394718 592692 394954
rect 592928 394718 592960 394954
rect -9036 394634 592960 394718
rect -9036 394398 -9004 394634
rect -8768 394398 -8684 394634
rect -8448 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592372 394634
rect 592608 394398 592692 394634
rect 592928 394398 592960 394634
rect -9036 394366 592960 394398
rect -9036 390454 592960 390486
rect -9036 390218 -8044 390454
rect -7808 390218 -7724 390454
rect -7488 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591412 390454
rect 591648 390218 591732 390454
rect 591968 390218 592960 390454
rect -9036 390134 592960 390218
rect -9036 389898 -8044 390134
rect -7808 389898 -7724 390134
rect -7488 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591412 390134
rect 591648 389898 591732 390134
rect 591968 389898 592960 390134
rect -9036 389866 592960 389898
rect -9036 385954 592960 385986
rect -9036 385718 -7084 385954
rect -6848 385718 -6764 385954
rect -6528 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590452 385954
rect 590688 385718 590772 385954
rect 591008 385718 592960 385954
rect -9036 385634 592960 385718
rect -9036 385398 -7084 385634
rect -6848 385398 -6764 385634
rect -6528 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590452 385634
rect 590688 385398 590772 385634
rect 591008 385398 592960 385634
rect -9036 385366 592960 385398
rect -9036 381454 592960 381486
rect -9036 381218 -6124 381454
rect -5888 381218 -5804 381454
rect -5568 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589492 381454
rect 589728 381218 589812 381454
rect 590048 381218 592960 381454
rect -9036 381134 592960 381218
rect -9036 380898 -6124 381134
rect -5888 380898 -5804 381134
rect -5568 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589492 381134
rect 589728 380898 589812 381134
rect 590048 380898 592960 381134
rect -9036 380866 592960 380898
rect -9036 376954 592960 376986
rect -9036 376718 -5164 376954
rect -4928 376718 -4844 376954
rect -4608 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588532 376954
rect 588768 376718 588852 376954
rect 589088 376718 592960 376954
rect -9036 376634 592960 376718
rect -9036 376398 -5164 376634
rect -4928 376398 -4844 376634
rect -4608 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588532 376634
rect 588768 376398 588852 376634
rect 589088 376398 592960 376634
rect -9036 376366 592960 376398
rect -9036 372454 592960 372486
rect -9036 372218 -4204 372454
rect -3968 372218 -3884 372454
rect -3648 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587572 372454
rect 587808 372218 587892 372454
rect 588128 372218 592960 372454
rect -9036 372134 592960 372218
rect -9036 371898 -4204 372134
rect -3968 371898 -3884 372134
rect -3648 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587572 372134
rect 587808 371898 587892 372134
rect 588128 371898 592960 372134
rect -9036 371866 592960 371898
rect -9036 367954 592960 367986
rect -9036 367718 -3244 367954
rect -3008 367718 -2924 367954
rect -2688 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586612 367954
rect 586848 367718 586932 367954
rect 587168 367718 592960 367954
rect -9036 367634 592960 367718
rect -9036 367398 -3244 367634
rect -3008 367398 -2924 367634
rect -2688 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586612 367634
rect 586848 367398 586932 367634
rect 587168 367398 592960 367634
rect -9036 367366 592960 367398
rect -9036 363454 592960 363486
rect -9036 363218 -2284 363454
rect -2048 363218 -1964 363454
rect -1728 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585652 363454
rect 585888 363218 585972 363454
rect 586208 363218 592960 363454
rect -9036 363134 592960 363218
rect -9036 362898 -2284 363134
rect -2048 362898 -1964 363134
rect -1728 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585652 363134
rect 585888 362898 585972 363134
rect 586208 362898 592960 363134
rect -9036 362866 592960 362898
rect -9036 358954 592960 358986
rect -9036 358718 -9004 358954
rect -8768 358718 -8684 358954
rect -8448 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592372 358954
rect 592608 358718 592692 358954
rect 592928 358718 592960 358954
rect -9036 358634 592960 358718
rect -9036 358398 -9004 358634
rect -8768 358398 -8684 358634
rect -8448 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592372 358634
rect 592608 358398 592692 358634
rect 592928 358398 592960 358634
rect -9036 358366 592960 358398
rect -9036 354454 592960 354486
rect -9036 354218 -8044 354454
rect -7808 354218 -7724 354454
rect -7488 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591412 354454
rect 591648 354218 591732 354454
rect 591968 354218 592960 354454
rect -9036 354134 592960 354218
rect -9036 353898 -8044 354134
rect -7808 353898 -7724 354134
rect -7488 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591412 354134
rect 591648 353898 591732 354134
rect 591968 353898 592960 354134
rect -9036 353866 592960 353898
rect -9036 349954 592960 349986
rect -9036 349718 -7084 349954
rect -6848 349718 -6764 349954
rect -6528 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590452 349954
rect 590688 349718 590772 349954
rect 591008 349718 592960 349954
rect -9036 349634 592960 349718
rect -9036 349398 -7084 349634
rect -6848 349398 -6764 349634
rect -6528 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590452 349634
rect 590688 349398 590772 349634
rect 591008 349398 592960 349634
rect -9036 349366 592960 349398
rect -9036 345454 592960 345486
rect -9036 345218 -6124 345454
rect -5888 345218 -5804 345454
rect -5568 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589492 345454
rect 589728 345218 589812 345454
rect 590048 345218 592960 345454
rect -9036 345134 592960 345218
rect -9036 344898 -6124 345134
rect -5888 344898 -5804 345134
rect -5568 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589492 345134
rect 589728 344898 589812 345134
rect 590048 344898 592960 345134
rect -9036 344866 592960 344898
rect -9036 340954 592960 340986
rect -9036 340718 -5164 340954
rect -4928 340718 -4844 340954
rect -4608 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588532 340954
rect 588768 340718 588852 340954
rect 589088 340718 592960 340954
rect -9036 340634 592960 340718
rect -9036 340398 -5164 340634
rect -4928 340398 -4844 340634
rect -4608 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588532 340634
rect 588768 340398 588852 340634
rect 589088 340398 592960 340634
rect -9036 340366 592960 340398
rect -9036 336454 592960 336486
rect -9036 336218 -4204 336454
rect -3968 336218 -3884 336454
rect -3648 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587572 336454
rect 587808 336218 587892 336454
rect 588128 336218 592960 336454
rect -9036 336134 592960 336218
rect -9036 335898 -4204 336134
rect -3968 335898 -3884 336134
rect -3648 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587572 336134
rect 587808 335898 587892 336134
rect 588128 335898 592960 336134
rect -9036 335866 592960 335898
rect -9036 331954 592960 331986
rect -9036 331718 -3244 331954
rect -3008 331718 -2924 331954
rect -2688 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586612 331954
rect 586848 331718 586932 331954
rect 587168 331718 592960 331954
rect -9036 331634 592960 331718
rect -9036 331398 -3244 331634
rect -3008 331398 -2924 331634
rect -2688 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586612 331634
rect 586848 331398 586932 331634
rect 587168 331398 592960 331634
rect -9036 331366 592960 331398
rect -9036 327454 592960 327486
rect -9036 327218 -2284 327454
rect -2048 327218 -1964 327454
rect -1728 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585652 327454
rect 585888 327218 585972 327454
rect 586208 327218 592960 327454
rect -9036 327134 592960 327218
rect -9036 326898 -2284 327134
rect -2048 326898 -1964 327134
rect -1728 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585652 327134
rect 585888 326898 585972 327134
rect 586208 326898 592960 327134
rect -9036 326866 592960 326898
rect -9036 322954 592960 322986
rect -9036 322718 -9004 322954
rect -8768 322718 -8684 322954
rect -8448 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592372 322954
rect 592608 322718 592692 322954
rect 592928 322718 592960 322954
rect -9036 322634 592960 322718
rect -9036 322398 -9004 322634
rect -8768 322398 -8684 322634
rect -8448 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592372 322634
rect 592608 322398 592692 322634
rect 592928 322398 592960 322634
rect -9036 322366 592960 322398
rect -9036 318454 592960 318486
rect -9036 318218 -8044 318454
rect -7808 318218 -7724 318454
rect -7488 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591412 318454
rect 591648 318218 591732 318454
rect 591968 318218 592960 318454
rect -9036 318134 592960 318218
rect -9036 317898 -8044 318134
rect -7808 317898 -7724 318134
rect -7488 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591412 318134
rect 591648 317898 591732 318134
rect 591968 317898 592960 318134
rect -9036 317866 592960 317898
rect -9036 313954 592960 313986
rect -9036 313718 -7084 313954
rect -6848 313718 -6764 313954
rect -6528 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590452 313954
rect 590688 313718 590772 313954
rect 591008 313718 592960 313954
rect -9036 313634 592960 313718
rect -9036 313398 -7084 313634
rect -6848 313398 -6764 313634
rect -6528 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590452 313634
rect 590688 313398 590772 313634
rect 591008 313398 592960 313634
rect -9036 313366 592960 313398
rect -9036 309454 592960 309486
rect -9036 309218 -6124 309454
rect -5888 309218 -5804 309454
rect -5568 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589492 309454
rect 589728 309218 589812 309454
rect 590048 309218 592960 309454
rect -9036 309134 592960 309218
rect -9036 308898 -6124 309134
rect -5888 308898 -5804 309134
rect -5568 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589492 309134
rect 589728 308898 589812 309134
rect 590048 308898 592960 309134
rect -9036 308866 592960 308898
rect -9036 304954 592960 304986
rect -9036 304718 -5164 304954
rect -4928 304718 -4844 304954
rect -4608 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588532 304954
rect 588768 304718 588852 304954
rect 589088 304718 592960 304954
rect -9036 304634 592960 304718
rect -9036 304398 -5164 304634
rect -4928 304398 -4844 304634
rect -4608 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588532 304634
rect 588768 304398 588852 304634
rect 589088 304398 592960 304634
rect -9036 304366 592960 304398
rect -9036 300454 592960 300486
rect -9036 300218 -4204 300454
rect -3968 300218 -3884 300454
rect -3648 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587572 300454
rect 587808 300218 587892 300454
rect 588128 300218 592960 300454
rect -9036 300134 592960 300218
rect -9036 299898 -4204 300134
rect -3968 299898 -3884 300134
rect -3648 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587572 300134
rect 587808 299898 587892 300134
rect 588128 299898 592960 300134
rect -9036 299866 592960 299898
rect -9036 295954 592960 295986
rect -9036 295718 -3244 295954
rect -3008 295718 -2924 295954
rect -2688 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586612 295954
rect 586848 295718 586932 295954
rect 587168 295718 592960 295954
rect -9036 295634 592960 295718
rect -9036 295398 -3244 295634
rect -3008 295398 -2924 295634
rect -2688 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586612 295634
rect 586848 295398 586932 295634
rect 587168 295398 592960 295634
rect -9036 295366 592960 295398
rect -9036 291454 592960 291486
rect -9036 291218 -2284 291454
rect -2048 291218 -1964 291454
rect -1728 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585652 291454
rect 585888 291218 585972 291454
rect 586208 291218 592960 291454
rect -9036 291134 592960 291218
rect -9036 290898 -2284 291134
rect -2048 290898 -1964 291134
rect -1728 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585652 291134
rect 585888 290898 585972 291134
rect 586208 290898 592960 291134
rect -9036 290866 592960 290898
rect -9036 286954 592960 286986
rect -9036 286718 -9004 286954
rect -8768 286718 -8684 286954
rect -8448 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592372 286954
rect 592608 286718 592692 286954
rect 592928 286718 592960 286954
rect -9036 286634 592960 286718
rect -9036 286398 -9004 286634
rect -8768 286398 -8684 286634
rect -8448 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592372 286634
rect 592608 286398 592692 286634
rect 592928 286398 592960 286634
rect -9036 286366 592960 286398
rect -9036 282454 592960 282486
rect -9036 282218 -8044 282454
rect -7808 282218 -7724 282454
rect -7488 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591412 282454
rect 591648 282218 591732 282454
rect 591968 282218 592960 282454
rect -9036 282134 592960 282218
rect -9036 281898 -8044 282134
rect -7808 281898 -7724 282134
rect -7488 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591412 282134
rect 591648 281898 591732 282134
rect 591968 281898 592960 282134
rect -9036 281866 592960 281898
rect -9036 277954 592960 277986
rect -9036 277718 -7084 277954
rect -6848 277718 -6764 277954
rect -6528 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590452 277954
rect 590688 277718 590772 277954
rect 591008 277718 592960 277954
rect -9036 277634 592960 277718
rect -9036 277398 -7084 277634
rect -6848 277398 -6764 277634
rect -6528 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590452 277634
rect 590688 277398 590772 277634
rect 591008 277398 592960 277634
rect -9036 277366 592960 277398
rect -9036 273454 592960 273486
rect -9036 273218 -6124 273454
rect -5888 273218 -5804 273454
rect -5568 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589492 273454
rect 589728 273218 589812 273454
rect 590048 273218 592960 273454
rect -9036 273134 592960 273218
rect -9036 272898 -6124 273134
rect -5888 272898 -5804 273134
rect -5568 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589492 273134
rect 589728 272898 589812 273134
rect 590048 272898 592960 273134
rect -9036 272866 592960 272898
rect -9036 268954 592960 268986
rect -9036 268718 -5164 268954
rect -4928 268718 -4844 268954
rect -4608 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588532 268954
rect 588768 268718 588852 268954
rect 589088 268718 592960 268954
rect -9036 268634 592960 268718
rect -9036 268398 -5164 268634
rect -4928 268398 -4844 268634
rect -4608 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588532 268634
rect 588768 268398 588852 268634
rect 589088 268398 592960 268634
rect -9036 268366 592960 268398
rect -9036 264454 592960 264486
rect -9036 264218 -4204 264454
rect -3968 264218 -3884 264454
rect -3648 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587572 264454
rect 587808 264218 587892 264454
rect 588128 264218 592960 264454
rect -9036 264134 592960 264218
rect -9036 263898 -4204 264134
rect -3968 263898 -3884 264134
rect -3648 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587572 264134
rect 587808 263898 587892 264134
rect 588128 263898 592960 264134
rect -9036 263866 592960 263898
rect -9036 259954 592960 259986
rect -9036 259718 -3244 259954
rect -3008 259718 -2924 259954
rect -2688 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586612 259954
rect 586848 259718 586932 259954
rect 587168 259718 592960 259954
rect -9036 259634 592960 259718
rect -9036 259398 -3244 259634
rect -3008 259398 -2924 259634
rect -2688 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586612 259634
rect 586848 259398 586932 259634
rect 587168 259398 592960 259634
rect -9036 259366 592960 259398
rect -9036 255454 592960 255486
rect -9036 255218 -2284 255454
rect -2048 255218 -1964 255454
rect -1728 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585652 255454
rect 585888 255218 585972 255454
rect 586208 255218 592960 255454
rect -9036 255134 592960 255218
rect -9036 254898 -2284 255134
rect -2048 254898 -1964 255134
rect -1728 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585652 255134
rect 585888 254898 585972 255134
rect 586208 254898 592960 255134
rect -9036 254866 592960 254898
rect -9036 250954 592960 250986
rect -9036 250718 -9004 250954
rect -8768 250718 -8684 250954
rect -8448 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592372 250954
rect 592608 250718 592692 250954
rect 592928 250718 592960 250954
rect -9036 250634 592960 250718
rect -9036 250398 -9004 250634
rect -8768 250398 -8684 250634
rect -8448 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592372 250634
rect 592608 250398 592692 250634
rect 592928 250398 592960 250634
rect -9036 250366 592960 250398
rect -9036 246454 592960 246486
rect -9036 246218 -8044 246454
rect -7808 246218 -7724 246454
rect -7488 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591412 246454
rect 591648 246218 591732 246454
rect 591968 246218 592960 246454
rect -9036 246134 592960 246218
rect -9036 245898 -8044 246134
rect -7808 245898 -7724 246134
rect -7488 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591412 246134
rect 591648 245898 591732 246134
rect 591968 245898 592960 246134
rect -9036 245866 592960 245898
rect -9036 241954 592960 241986
rect -9036 241718 -7084 241954
rect -6848 241718 -6764 241954
rect -6528 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590452 241954
rect 590688 241718 590772 241954
rect 591008 241718 592960 241954
rect -9036 241634 592960 241718
rect -9036 241398 -7084 241634
rect -6848 241398 -6764 241634
rect -6528 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590452 241634
rect 590688 241398 590772 241634
rect 591008 241398 592960 241634
rect -9036 241366 592960 241398
rect -9036 237454 592960 237486
rect -9036 237218 -6124 237454
rect -5888 237218 -5804 237454
rect -5568 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589492 237454
rect 589728 237218 589812 237454
rect 590048 237218 592960 237454
rect -9036 237134 592960 237218
rect -9036 236898 -6124 237134
rect -5888 236898 -5804 237134
rect -5568 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589492 237134
rect 589728 236898 589812 237134
rect 590048 236898 592960 237134
rect -9036 236866 592960 236898
rect -9036 232954 592960 232986
rect -9036 232718 -5164 232954
rect -4928 232718 -4844 232954
rect -4608 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588532 232954
rect 588768 232718 588852 232954
rect 589088 232718 592960 232954
rect -9036 232634 592960 232718
rect -9036 232398 -5164 232634
rect -4928 232398 -4844 232634
rect -4608 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588532 232634
rect 588768 232398 588852 232634
rect 589088 232398 592960 232634
rect -9036 232366 592960 232398
rect -9036 228454 592960 228486
rect -9036 228218 -4204 228454
rect -3968 228218 -3884 228454
rect -3648 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587572 228454
rect 587808 228218 587892 228454
rect 588128 228218 592960 228454
rect -9036 228134 592960 228218
rect -9036 227898 -4204 228134
rect -3968 227898 -3884 228134
rect -3648 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587572 228134
rect 587808 227898 587892 228134
rect 588128 227898 592960 228134
rect -9036 227866 592960 227898
rect -9036 223954 592960 223986
rect -9036 223718 -3244 223954
rect -3008 223718 -2924 223954
rect -2688 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586612 223954
rect 586848 223718 586932 223954
rect 587168 223718 592960 223954
rect -9036 223634 592960 223718
rect -9036 223398 -3244 223634
rect -3008 223398 -2924 223634
rect -2688 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586612 223634
rect 586848 223398 586932 223634
rect 587168 223398 592960 223634
rect -9036 223366 592960 223398
rect -9036 219454 592960 219486
rect -9036 219218 -2284 219454
rect -2048 219218 -1964 219454
rect -1728 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585652 219454
rect 585888 219218 585972 219454
rect 586208 219218 592960 219454
rect -9036 219134 592960 219218
rect -9036 218898 -2284 219134
rect -2048 218898 -1964 219134
rect -1728 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585652 219134
rect 585888 218898 585972 219134
rect 586208 218898 592960 219134
rect -9036 218866 592960 218898
rect -9036 214954 592960 214986
rect -9036 214718 -9004 214954
rect -8768 214718 -8684 214954
rect -8448 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592372 214954
rect 592608 214718 592692 214954
rect 592928 214718 592960 214954
rect -9036 214634 592960 214718
rect -9036 214398 -9004 214634
rect -8768 214398 -8684 214634
rect -8448 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592372 214634
rect 592608 214398 592692 214634
rect 592928 214398 592960 214634
rect -9036 214366 592960 214398
rect -9036 210454 592960 210486
rect -9036 210218 -8044 210454
rect -7808 210218 -7724 210454
rect -7488 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591412 210454
rect 591648 210218 591732 210454
rect 591968 210218 592960 210454
rect -9036 210134 592960 210218
rect -9036 209898 -8044 210134
rect -7808 209898 -7724 210134
rect -7488 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591412 210134
rect 591648 209898 591732 210134
rect 591968 209898 592960 210134
rect -9036 209866 592960 209898
rect -9036 205954 592960 205986
rect -9036 205718 -7084 205954
rect -6848 205718 -6764 205954
rect -6528 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590452 205954
rect 590688 205718 590772 205954
rect 591008 205718 592960 205954
rect -9036 205634 592960 205718
rect -9036 205398 -7084 205634
rect -6848 205398 -6764 205634
rect -6528 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590452 205634
rect 590688 205398 590772 205634
rect 591008 205398 592960 205634
rect -9036 205366 592960 205398
rect -9036 201454 592960 201486
rect -9036 201218 -6124 201454
rect -5888 201218 -5804 201454
rect -5568 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589492 201454
rect 589728 201218 589812 201454
rect 590048 201218 592960 201454
rect -9036 201134 592960 201218
rect -9036 200898 -6124 201134
rect -5888 200898 -5804 201134
rect -5568 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589492 201134
rect 589728 200898 589812 201134
rect 590048 200898 592960 201134
rect -9036 200866 592960 200898
rect -9036 196954 592960 196986
rect -9036 196718 -5164 196954
rect -4928 196718 -4844 196954
rect -4608 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588532 196954
rect 588768 196718 588852 196954
rect 589088 196718 592960 196954
rect -9036 196634 592960 196718
rect -9036 196398 -5164 196634
rect -4928 196398 -4844 196634
rect -4608 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588532 196634
rect 588768 196398 588852 196634
rect 589088 196398 592960 196634
rect -9036 196366 592960 196398
rect -9036 192454 592960 192486
rect -9036 192218 -4204 192454
rect -3968 192218 -3884 192454
rect -3648 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587572 192454
rect 587808 192218 587892 192454
rect 588128 192218 592960 192454
rect -9036 192134 592960 192218
rect -9036 191898 -4204 192134
rect -3968 191898 -3884 192134
rect -3648 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587572 192134
rect 587808 191898 587892 192134
rect 588128 191898 592960 192134
rect -9036 191866 592960 191898
rect -9036 187954 592960 187986
rect -9036 187718 -3244 187954
rect -3008 187718 -2924 187954
rect -2688 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586612 187954
rect 586848 187718 586932 187954
rect 587168 187718 592960 187954
rect -9036 187634 592960 187718
rect -9036 187398 -3244 187634
rect -3008 187398 -2924 187634
rect -2688 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586612 187634
rect 586848 187398 586932 187634
rect 587168 187398 592960 187634
rect -9036 187366 592960 187398
rect -9036 183454 592960 183486
rect -9036 183218 -2284 183454
rect -2048 183218 -1964 183454
rect -1728 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585652 183454
rect 585888 183218 585972 183454
rect 586208 183218 592960 183454
rect -9036 183134 592960 183218
rect -9036 182898 -2284 183134
rect -2048 182898 -1964 183134
rect -1728 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585652 183134
rect 585888 182898 585972 183134
rect 586208 182898 592960 183134
rect -9036 182866 592960 182898
rect -9036 178954 592960 178986
rect -9036 178718 -9004 178954
rect -8768 178718 -8684 178954
rect -8448 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592372 178954
rect 592608 178718 592692 178954
rect 592928 178718 592960 178954
rect -9036 178634 592960 178718
rect -9036 178398 -9004 178634
rect -8768 178398 -8684 178634
rect -8448 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592372 178634
rect 592608 178398 592692 178634
rect 592928 178398 592960 178634
rect -9036 178366 592960 178398
rect -9036 174454 592960 174486
rect -9036 174218 -8044 174454
rect -7808 174218 -7724 174454
rect -7488 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591412 174454
rect 591648 174218 591732 174454
rect 591968 174218 592960 174454
rect -9036 174134 592960 174218
rect -9036 173898 -8044 174134
rect -7808 173898 -7724 174134
rect -7488 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591412 174134
rect 591648 173898 591732 174134
rect 591968 173898 592960 174134
rect -9036 173866 592960 173898
rect -9036 169954 592960 169986
rect -9036 169718 -7084 169954
rect -6848 169718 -6764 169954
rect -6528 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590452 169954
rect 590688 169718 590772 169954
rect 591008 169718 592960 169954
rect -9036 169634 592960 169718
rect -9036 169398 -7084 169634
rect -6848 169398 -6764 169634
rect -6528 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590452 169634
rect 590688 169398 590772 169634
rect 591008 169398 592960 169634
rect -9036 169366 592960 169398
rect -9036 165454 592960 165486
rect -9036 165218 -6124 165454
rect -5888 165218 -5804 165454
rect -5568 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589492 165454
rect 589728 165218 589812 165454
rect 590048 165218 592960 165454
rect -9036 165134 592960 165218
rect -9036 164898 -6124 165134
rect -5888 164898 -5804 165134
rect -5568 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589492 165134
rect 589728 164898 589812 165134
rect 590048 164898 592960 165134
rect -9036 164866 592960 164898
rect -9036 160954 592960 160986
rect -9036 160718 -5164 160954
rect -4928 160718 -4844 160954
rect -4608 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588532 160954
rect 588768 160718 588852 160954
rect 589088 160718 592960 160954
rect -9036 160634 592960 160718
rect -9036 160398 -5164 160634
rect -4928 160398 -4844 160634
rect -4608 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588532 160634
rect 588768 160398 588852 160634
rect 589088 160398 592960 160634
rect -9036 160366 592960 160398
rect -9036 156454 592960 156486
rect -9036 156218 -4204 156454
rect -3968 156218 -3884 156454
rect -3648 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587572 156454
rect 587808 156218 587892 156454
rect 588128 156218 592960 156454
rect -9036 156134 592960 156218
rect -9036 155898 -4204 156134
rect -3968 155898 -3884 156134
rect -3648 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587572 156134
rect 587808 155898 587892 156134
rect 588128 155898 592960 156134
rect -9036 155866 592960 155898
rect -9036 151954 592960 151986
rect -9036 151718 -3244 151954
rect -3008 151718 -2924 151954
rect -2688 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586612 151954
rect 586848 151718 586932 151954
rect 587168 151718 592960 151954
rect -9036 151634 592960 151718
rect -9036 151398 -3244 151634
rect -3008 151398 -2924 151634
rect -2688 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586612 151634
rect 586848 151398 586932 151634
rect 587168 151398 592960 151634
rect -9036 151366 592960 151398
rect -9036 147454 592960 147486
rect -9036 147218 -2284 147454
rect -2048 147218 -1964 147454
rect -1728 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147239 145826 147454
rect 74382 147218 84250 147239
rect -9036 147134 84250 147218
rect -9036 146898 -2284 147134
rect -2048 146898 -1964 147134
rect -1728 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 147003 84250 147134
rect 84486 147003 114970 147239
rect 115206 147218 145826 147239
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585652 147454
rect 585888 147218 585972 147454
rect 586208 147218 592960 147454
rect 115206 147134 592960 147218
rect 115206 147003 145826 147134
rect 74382 146898 145826 147003
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585652 147134
rect 585888 146898 585972 147134
rect 586208 146898 592960 147134
rect -9036 146866 592960 146898
rect -9036 142954 592960 142986
rect -9036 142718 -9004 142954
rect -8768 142718 -8684 142954
rect -8448 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592372 142954
rect 592608 142718 592692 142954
rect 592928 142718 592960 142954
rect -9036 142634 592960 142718
rect -9036 142398 -9004 142634
rect -8768 142398 -8684 142634
rect -8448 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592372 142634
rect 592608 142398 592692 142634
rect 592928 142398 592960 142634
rect -9036 142366 592960 142398
rect -9036 138454 592960 138486
rect -9036 138218 -8044 138454
rect -7808 138218 -7724 138454
rect -7488 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591412 138454
rect 591648 138218 591732 138454
rect 591968 138218 592960 138454
rect -9036 138134 592960 138218
rect -9036 137898 -8044 138134
rect -7808 137898 -7724 138134
rect -7488 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591412 138134
rect 591648 137898 591732 138134
rect 591968 137898 592960 138134
rect -9036 137866 592960 137898
rect -9036 133954 592960 133986
rect -9036 133718 -7084 133954
rect -6848 133718 -6764 133954
rect -6528 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590452 133954
rect 590688 133718 590772 133954
rect 591008 133718 592960 133954
rect -9036 133634 592960 133718
rect -9036 133398 -7084 133634
rect -6848 133398 -6764 133634
rect -6528 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590452 133634
rect 590688 133398 590772 133634
rect 591008 133398 592960 133634
rect -9036 133366 592960 133398
rect -9036 129454 592960 129486
rect -9036 129218 -6124 129454
rect -5888 129218 -5804 129454
rect -5568 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589492 129454
rect 589728 129218 589812 129454
rect 590048 129218 592960 129454
rect -9036 129134 592960 129218
rect -9036 128898 -6124 129134
rect -5888 128898 -5804 129134
rect -5568 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589492 129134
rect 589728 128898 589812 129134
rect 590048 128898 592960 129134
rect -9036 128866 592960 128898
rect -9036 124954 592960 124986
rect -9036 124718 -5164 124954
rect -4928 124718 -4844 124954
rect -4608 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588532 124954
rect 588768 124718 588852 124954
rect 589088 124718 592960 124954
rect -9036 124634 592960 124718
rect -9036 124398 -5164 124634
rect -4928 124398 -4844 124634
rect -4608 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588532 124634
rect 588768 124398 588852 124634
rect 589088 124398 592960 124634
rect -9036 124366 592960 124398
rect -9036 120454 592960 120486
rect -9036 120218 -4204 120454
rect -3968 120218 -3884 120454
rect -3648 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587572 120454
rect 587808 120218 587892 120454
rect 588128 120218 592960 120454
rect -9036 120134 592960 120218
rect -9036 119898 -4204 120134
rect -3968 119898 -3884 120134
rect -3648 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587572 120134
rect 587808 119898 587892 120134
rect 588128 119898 592960 120134
rect -9036 119866 592960 119898
rect -9036 115954 592960 115986
rect -9036 115718 -3244 115954
rect -3008 115718 -2924 115954
rect -2688 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 99610 115954
rect 99846 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586612 115954
rect 586848 115718 586932 115954
rect 587168 115718 592960 115954
rect -9036 115634 592960 115718
rect -9036 115398 -3244 115634
rect -3008 115398 -2924 115634
rect -2688 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 99610 115634
rect 99846 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586612 115634
rect 586848 115398 586932 115634
rect 587168 115398 592960 115634
rect -9036 115366 592960 115398
rect -9036 111454 592960 111486
rect -9036 111218 -2284 111454
rect -2048 111218 -1964 111454
rect -1728 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 84250 111454
rect 84486 111218 114970 111454
rect 115206 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585652 111454
rect 585888 111218 585972 111454
rect 586208 111218 592960 111454
rect -9036 111134 592960 111218
rect -9036 110898 -2284 111134
rect -2048 110898 -1964 111134
rect -1728 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 84250 111134
rect 84486 110898 114970 111134
rect 115206 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585652 111134
rect 585888 110898 585972 111134
rect 586208 110898 592960 111134
rect -9036 110866 592960 110898
rect -9036 106954 592960 106986
rect -9036 106718 -9004 106954
rect -8768 106718 -8684 106954
rect -8448 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592372 106954
rect 592608 106718 592692 106954
rect 592928 106718 592960 106954
rect -9036 106634 592960 106718
rect -9036 106398 -9004 106634
rect -8768 106398 -8684 106634
rect -8448 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592372 106634
rect 592608 106398 592692 106634
rect 592928 106398 592960 106634
rect -9036 106366 592960 106398
rect -9036 102454 592960 102486
rect -9036 102218 -8044 102454
rect -7808 102218 -7724 102454
rect -7488 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591412 102454
rect 591648 102218 591732 102454
rect 591968 102218 592960 102454
rect -9036 102134 592960 102218
rect -9036 101898 -8044 102134
rect -7808 101898 -7724 102134
rect -7488 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591412 102134
rect 591648 101898 591732 102134
rect 591968 101898 592960 102134
rect -9036 101866 592960 101898
rect -9036 97954 592960 97986
rect -9036 97718 -7084 97954
rect -6848 97718 -6764 97954
rect -6528 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590452 97954
rect 590688 97718 590772 97954
rect 591008 97718 592960 97954
rect -9036 97634 592960 97718
rect -9036 97398 -7084 97634
rect -6848 97398 -6764 97634
rect -6528 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590452 97634
rect 590688 97398 590772 97634
rect 591008 97398 592960 97634
rect -9036 97366 592960 97398
rect -9036 93454 592960 93486
rect -9036 93218 -6124 93454
rect -5888 93218 -5804 93454
rect -5568 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589492 93454
rect 589728 93218 589812 93454
rect 590048 93218 592960 93454
rect -9036 93134 592960 93218
rect -9036 92898 -6124 93134
rect -5888 92898 -5804 93134
rect -5568 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589492 93134
rect 589728 92898 589812 93134
rect 590048 92898 592960 93134
rect -9036 92866 592960 92898
rect -9036 88954 592960 88986
rect -9036 88718 -5164 88954
rect -4928 88718 -4844 88954
rect -4608 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588532 88954
rect 588768 88718 588852 88954
rect 589088 88718 592960 88954
rect -9036 88634 592960 88718
rect -9036 88398 -5164 88634
rect -4928 88398 -4844 88634
rect -4608 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588532 88634
rect 588768 88398 588852 88634
rect 589088 88398 592960 88634
rect -9036 88366 592960 88398
rect -9036 84454 592960 84486
rect -9036 84218 -4204 84454
rect -3968 84218 -3884 84454
rect -3648 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587572 84454
rect 587808 84218 587892 84454
rect 588128 84218 592960 84454
rect -9036 84134 592960 84218
rect -9036 83898 -4204 84134
rect -3968 83898 -3884 84134
rect -3648 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587572 84134
rect 587808 83898 587892 84134
rect 588128 83898 592960 84134
rect -9036 83866 592960 83898
rect -9036 79954 592960 79986
rect -9036 79718 -3244 79954
rect -3008 79718 -2924 79954
rect -2688 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586612 79954
rect 586848 79718 586932 79954
rect 587168 79718 592960 79954
rect -9036 79634 592960 79718
rect -9036 79398 -3244 79634
rect -3008 79398 -2924 79634
rect -2688 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586612 79634
rect 586848 79398 586932 79634
rect 587168 79398 592960 79634
rect -9036 79366 592960 79398
rect -9036 75454 592960 75486
rect -9036 75218 -2284 75454
rect -2048 75218 -1964 75454
rect -1728 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585652 75454
rect 585888 75218 585972 75454
rect 586208 75218 592960 75454
rect -9036 75134 592960 75218
rect -9036 74898 -2284 75134
rect -2048 74898 -1964 75134
rect -1728 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585652 75134
rect 585888 74898 585972 75134
rect 586208 74898 592960 75134
rect -9036 74866 592960 74898
rect -9036 70954 592960 70986
rect -9036 70718 -9004 70954
rect -8768 70718 -8684 70954
rect -8448 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592372 70954
rect 592608 70718 592692 70954
rect 592928 70718 592960 70954
rect -9036 70634 592960 70718
rect -9036 70398 -9004 70634
rect -8768 70398 -8684 70634
rect -8448 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592372 70634
rect 592608 70398 592692 70634
rect 592928 70398 592960 70634
rect -9036 70366 592960 70398
rect -9036 66454 592960 66486
rect -9036 66218 -8044 66454
rect -7808 66218 -7724 66454
rect -7488 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591412 66454
rect 591648 66218 591732 66454
rect 591968 66218 592960 66454
rect -9036 66134 592960 66218
rect -9036 65898 -8044 66134
rect -7808 65898 -7724 66134
rect -7488 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591412 66134
rect 591648 65898 591732 66134
rect 591968 65898 592960 66134
rect -9036 65866 592960 65898
rect -9036 61954 592960 61986
rect -9036 61718 -7084 61954
rect -6848 61718 -6764 61954
rect -6528 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590452 61954
rect 590688 61718 590772 61954
rect 591008 61718 592960 61954
rect -9036 61634 592960 61718
rect -9036 61398 -7084 61634
rect -6848 61398 -6764 61634
rect -6528 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590452 61634
rect 590688 61398 590772 61634
rect 591008 61398 592960 61634
rect -9036 61366 592960 61398
rect -9036 57454 592960 57486
rect -9036 57218 -6124 57454
rect -5888 57218 -5804 57454
rect -5568 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589492 57454
rect 589728 57218 589812 57454
rect 590048 57218 592960 57454
rect -9036 57134 592960 57218
rect -9036 56898 -6124 57134
rect -5888 56898 -5804 57134
rect -5568 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589492 57134
rect 589728 56898 589812 57134
rect 590048 56898 592960 57134
rect -9036 56866 592960 56898
rect -9036 52954 592960 52986
rect -9036 52718 -5164 52954
rect -4928 52718 -4844 52954
rect -4608 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588532 52954
rect 588768 52718 588852 52954
rect 589088 52718 592960 52954
rect -9036 52634 592960 52718
rect -9036 52398 -5164 52634
rect -4928 52398 -4844 52634
rect -4608 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588532 52634
rect 588768 52398 588852 52634
rect 589088 52398 592960 52634
rect -9036 52366 592960 52398
rect -9036 48454 592960 48486
rect -9036 48218 -4204 48454
rect -3968 48218 -3884 48454
rect -3648 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587572 48454
rect 587808 48218 587892 48454
rect 588128 48218 592960 48454
rect -9036 48134 592960 48218
rect -9036 47898 -4204 48134
rect -3968 47898 -3884 48134
rect -3648 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587572 48134
rect 587808 47898 587892 48134
rect 588128 47898 592960 48134
rect -9036 47866 592960 47898
rect -9036 43954 592960 43986
rect -9036 43718 -3244 43954
rect -3008 43718 -2924 43954
rect -2688 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586612 43954
rect 586848 43718 586932 43954
rect 587168 43718 592960 43954
rect -9036 43634 592960 43718
rect -9036 43398 -3244 43634
rect -3008 43398 -2924 43634
rect -2688 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586612 43634
rect 586848 43398 586932 43634
rect 587168 43398 592960 43634
rect -9036 43366 592960 43398
rect -9036 39454 592960 39486
rect -9036 39218 -2284 39454
rect -2048 39218 -1964 39454
rect -1728 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585652 39454
rect 585888 39218 585972 39454
rect 586208 39218 592960 39454
rect -9036 39134 592960 39218
rect -9036 38898 -2284 39134
rect -2048 38898 -1964 39134
rect -1728 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585652 39134
rect 585888 38898 585972 39134
rect 586208 38898 592960 39134
rect -9036 38866 592960 38898
rect -9036 34954 592960 34986
rect -9036 34718 -9004 34954
rect -8768 34718 -8684 34954
rect -8448 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592372 34954
rect 592608 34718 592692 34954
rect 592928 34718 592960 34954
rect -9036 34634 592960 34718
rect -9036 34398 -9004 34634
rect -8768 34398 -8684 34634
rect -8448 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592372 34634
rect 592608 34398 592692 34634
rect 592928 34398 592960 34634
rect -9036 34366 592960 34398
rect -9036 30454 592960 30486
rect -9036 30218 -8044 30454
rect -7808 30218 -7724 30454
rect -7488 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591412 30454
rect 591648 30218 591732 30454
rect 591968 30218 592960 30454
rect -9036 30134 592960 30218
rect -9036 29898 -8044 30134
rect -7808 29898 -7724 30134
rect -7488 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591412 30134
rect 591648 29898 591732 30134
rect 591968 29898 592960 30134
rect -9036 29866 592960 29898
rect -9036 25954 592960 25986
rect -9036 25718 -7084 25954
rect -6848 25718 -6764 25954
rect -6528 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590452 25954
rect 590688 25718 590772 25954
rect 591008 25718 592960 25954
rect -9036 25634 592960 25718
rect -9036 25398 -7084 25634
rect -6848 25398 -6764 25634
rect -6528 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590452 25634
rect 590688 25398 590772 25634
rect 591008 25398 592960 25634
rect -9036 25366 592960 25398
rect -9036 21454 592960 21486
rect -9036 21218 -6124 21454
rect -5888 21218 -5804 21454
rect -5568 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589492 21454
rect 589728 21218 589812 21454
rect 590048 21218 592960 21454
rect -9036 21134 592960 21218
rect -9036 20898 -6124 21134
rect -5888 20898 -5804 21134
rect -5568 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589492 21134
rect 589728 20898 589812 21134
rect 590048 20898 592960 21134
rect -9036 20866 592960 20898
rect -9036 16954 592960 16986
rect -9036 16718 -5164 16954
rect -4928 16718 -4844 16954
rect -4608 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588532 16954
rect 588768 16718 588852 16954
rect 589088 16718 592960 16954
rect -9036 16634 592960 16718
rect -9036 16398 -5164 16634
rect -4928 16398 -4844 16634
rect -4608 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588532 16634
rect 588768 16398 588852 16634
rect 589088 16398 592960 16634
rect -9036 16366 592960 16398
rect -9036 12454 592960 12486
rect -9036 12218 -4204 12454
rect -3968 12218 -3884 12454
rect -3648 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587572 12454
rect 587808 12218 587892 12454
rect 588128 12218 592960 12454
rect -9036 12134 592960 12218
rect -9036 11898 -4204 12134
rect -3968 11898 -3884 12134
rect -3648 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587572 12134
rect 587808 11898 587892 12134
rect 588128 11898 592960 12134
rect -9036 11866 592960 11898
rect -9036 7954 592960 7986
rect -9036 7718 -3244 7954
rect -3008 7718 -2924 7954
rect -2688 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586612 7954
rect 586848 7718 586932 7954
rect 587168 7718 592960 7954
rect -9036 7634 592960 7718
rect -9036 7398 -3244 7634
rect -3008 7398 -2924 7634
rect -2688 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586612 7634
rect 586848 7398 586932 7634
rect 587168 7398 592960 7634
rect -9036 7366 592960 7398
rect -9036 3454 592960 3486
rect -9036 3218 -2284 3454
rect -2048 3218 -1964 3454
rect -1728 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585652 3454
rect 585888 3218 585972 3454
rect 586208 3218 592960 3454
rect -9036 3134 592960 3218
rect -9036 2898 -2284 3134
rect -2048 2898 -1964 3134
rect -1728 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585652 3134
rect 585888 2898 585972 3134
rect 586208 2898 592960 3134
rect -9036 2866 592960 2898
rect -2316 -656 586240 -624
rect -2316 -892 -2284 -656
rect -2048 -892 -1964 -656
rect -1728 -892 1826 -656
rect 2062 -892 2146 -656
rect 2382 -892 37826 -656
rect 38062 -892 38146 -656
rect 38382 -892 73826 -656
rect 74062 -892 74146 -656
rect 74382 -892 109826 -656
rect 110062 -892 110146 -656
rect 110382 -892 145826 -656
rect 146062 -892 146146 -656
rect 146382 -892 181826 -656
rect 182062 -892 182146 -656
rect 182382 -892 217826 -656
rect 218062 -892 218146 -656
rect 218382 -892 253826 -656
rect 254062 -892 254146 -656
rect 254382 -892 289826 -656
rect 290062 -892 290146 -656
rect 290382 -892 325826 -656
rect 326062 -892 326146 -656
rect 326382 -892 361826 -656
rect 362062 -892 362146 -656
rect 362382 -892 397826 -656
rect 398062 -892 398146 -656
rect 398382 -892 433826 -656
rect 434062 -892 434146 -656
rect 434382 -892 469826 -656
rect 470062 -892 470146 -656
rect 470382 -892 505826 -656
rect 506062 -892 506146 -656
rect 506382 -892 541826 -656
rect 542062 -892 542146 -656
rect 542382 -892 577826 -656
rect 578062 -892 578146 -656
rect 578382 -892 585652 -656
rect 585888 -892 585972 -656
rect 586208 -892 586240 -656
rect -2316 -976 586240 -892
rect -2316 -1212 -2284 -976
rect -2048 -1212 -1964 -976
rect -1728 -1212 1826 -976
rect 2062 -1212 2146 -976
rect 2382 -1212 37826 -976
rect 38062 -1212 38146 -976
rect 38382 -1212 73826 -976
rect 74062 -1212 74146 -976
rect 74382 -1212 109826 -976
rect 110062 -1212 110146 -976
rect 110382 -1212 145826 -976
rect 146062 -1212 146146 -976
rect 146382 -1212 181826 -976
rect 182062 -1212 182146 -976
rect 182382 -1212 217826 -976
rect 218062 -1212 218146 -976
rect 218382 -1212 253826 -976
rect 254062 -1212 254146 -976
rect 254382 -1212 289826 -976
rect 290062 -1212 290146 -976
rect 290382 -1212 325826 -976
rect 326062 -1212 326146 -976
rect 326382 -1212 361826 -976
rect 362062 -1212 362146 -976
rect 362382 -1212 397826 -976
rect 398062 -1212 398146 -976
rect 398382 -1212 433826 -976
rect 434062 -1212 434146 -976
rect 434382 -1212 469826 -976
rect 470062 -1212 470146 -976
rect 470382 -1212 505826 -976
rect 506062 -1212 506146 -976
rect 506382 -1212 541826 -976
rect 542062 -1212 542146 -976
rect 542382 -1212 577826 -976
rect 578062 -1212 578146 -976
rect 578382 -1212 585652 -976
rect 585888 -1212 585972 -976
rect 586208 -1212 586240 -976
rect -2316 -1244 586240 -1212
rect -3276 -1616 587200 -1584
rect -3276 -1852 -3244 -1616
rect -3008 -1852 -2924 -1616
rect -2688 -1852 6326 -1616
rect 6562 -1852 6646 -1616
rect 6882 -1852 42326 -1616
rect 42562 -1852 42646 -1616
rect 42882 -1852 78326 -1616
rect 78562 -1852 78646 -1616
rect 78882 -1852 114326 -1616
rect 114562 -1852 114646 -1616
rect 114882 -1852 150326 -1616
rect 150562 -1852 150646 -1616
rect 150882 -1852 186326 -1616
rect 186562 -1852 186646 -1616
rect 186882 -1852 222326 -1616
rect 222562 -1852 222646 -1616
rect 222882 -1852 258326 -1616
rect 258562 -1852 258646 -1616
rect 258882 -1852 294326 -1616
rect 294562 -1852 294646 -1616
rect 294882 -1852 330326 -1616
rect 330562 -1852 330646 -1616
rect 330882 -1852 366326 -1616
rect 366562 -1852 366646 -1616
rect 366882 -1852 402326 -1616
rect 402562 -1852 402646 -1616
rect 402882 -1852 438326 -1616
rect 438562 -1852 438646 -1616
rect 438882 -1852 474326 -1616
rect 474562 -1852 474646 -1616
rect 474882 -1852 510326 -1616
rect 510562 -1852 510646 -1616
rect 510882 -1852 546326 -1616
rect 546562 -1852 546646 -1616
rect 546882 -1852 582326 -1616
rect 582562 -1852 582646 -1616
rect 582882 -1852 586612 -1616
rect 586848 -1852 586932 -1616
rect 587168 -1852 587200 -1616
rect -3276 -1936 587200 -1852
rect -3276 -2172 -3244 -1936
rect -3008 -2172 -2924 -1936
rect -2688 -2172 6326 -1936
rect 6562 -2172 6646 -1936
rect 6882 -2172 42326 -1936
rect 42562 -2172 42646 -1936
rect 42882 -2172 78326 -1936
rect 78562 -2172 78646 -1936
rect 78882 -2172 114326 -1936
rect 114562 -2172 114646 -1936
rect 114882 -2172 150326 -1936
rect 150562 -2172 150646 -1936
rect 150882 -2172 186326 -1936
rect 186562 -2172 186646 -1936
rect 186882 -2172 222326 -1936
rect 222562 -2172 222646 -1936
rect 222882 -2172 258326 -1936
rect 258562 -2172 258646 -1936
rect 258882 -2172 294326 -1936
rect 294562 -2172 294646 -1936
rect 294882 -2172 330326 -1936
rect 330562 -2172 330646 -1936
rect 330882 -2172 366326 -1936
rect 366562 -2172 366646 -1936
rect 366882 -2172 402326 -1936
rect 402562 -2172 402646 -1936
rect 402882 -2172 438326 -1936
rect 438562 -2172 438646 -1936
rect 438882 -2172 474326 -1936
rect 474562 -2172 474646 -1936
rect 474882 -2172 510326 -1936
rect 510562 -2172 510646 -1936
rect 510882 -2172 546326 -1936
rect 546562 -2172 546646 -1936
rect 546882 -2172 582326 -1936
rect 582562 -2172 582646 -1936
rect 582882 -2172 586612 -1936
rect 586848 -2172 586932 -1936
rect 587168 -2172 587200 -1936
rect -3276 -2204 587200 -2172
rect -4236 -2576 588160 -2544
rect -4236 -2812 -4204 -2576
rect -3968 -2812 -3884 -2576
rect -3648 -2812 10826 -2576
rect 11062 -2812 11146 -2576
rect 11382 -2812 46826 -2576
rect 47062 -2812 47146 -2576
rect 47382 -2812 82826 -2576
rect 83062 -2812 83146 -2576
rect 83382 -2812 118826 -2576
rect 119062 -2812 119146 -2576
rect 119382 -2812 154826 -2576
rect 155062 -2812 155146 -2576
rect 155382 -2812 190826 -2576
rect 191062 -2812 191146 -2576
rect 191382 -2812 226826 -2576
rect 227062 -2812 227146 -2576
rect 227382 -2812 262826 -2576
rect 263062 -2812 263146 -2576
rect 263382 -2812 298826 -2576
rect 299062 -2812 299146 -2576
rect 299382 -2812 334826 -2576
rect 335062 -2812 335146 -2576
rect 335382 -2812 370826 -2576
rect 371062 -2812 371146 -2576
rect 371382 -2812 406826 -2576
rect 407062 -2812 407146 -2576
rect 407382 -2812 442826 -2576
rect 443062 -2812 443146 -2576
rect 443382 -2812 478826 -2576
rect 479062 -2812 479146 -2576
rect 479382 -2812 514826 -2576
rect 515062 -2812 515146 -2576
rect 515382 -2812 550826 -2576
rect 551062 -2812 551146 -2576
rect 551382 -2812 587572 -2576
rect 587808 -2812 587892 -2576
rect 588128 -2812 588160 -2576
rect -4236 -2896 588160 -2812
rect -4236 -3132 -4204 -2896
rect -3968 -3132 -3884 -2896
rect -3648 -3132 10826 -2896
rect 11062 -3132 11146 -2896
rect 11382 -3132 46826 -2896
rect 47062 -3132 47146 -2896
rect 47382 -3132 82826 -2896
rect 83062 -3132 83146 -2896
rect 83382 -3132 118826 -2896
rect 119062 -3132 119146 -2896
rect 119382 -3132 154826 -2896
rect 155062 -3132 155146 -2896
rect 155382 -3132 190826 -2896
rect 191062 -3132 191146 -2896
rect 191382 -3132 226826 -2896
rect 227062 -3132 227146 -2896
rect 227382 -3132 262826 -2896
rect 263062 -3132 263146 -2896
rect 263382 -3132 298826 -2896
rect 299062 -3132 299146 -2896
rect 299382 -3132 334826 -2896
rect 335062 -3132 335146 -2896
rect 335382 -3132 370826 -2896
rect 371062 -3132 371146 -2896
rect 371382 -3132 406826 -2896
rect 407062 -3132 407146 -2896
rect 407382 -3132 442826 -2896
rect 443062 -3132 443146 -2896
rect 443382 -3132 478826 -2896
rect 479062 -3132 479146 -2896
rect 479382 -3132 514826 -2896
rect 515062 -3132 515146 -2896
rect 515382 -3132 550826 -2896
rect 551062 -3132 551146 -2896
rect 551382 -3132 587572 -2896
rect 587808 -3132 587892 -2896
rect 588128 -3132 588160 -2896
rect -4236 -3164 588160 -3132
rect -5196 -3536 589120 -3504
rect -5196 -3772 -5164 -3536
rect -4928 -3772 -4844 -3536
rect -4608 -3772 15326 -3536
rect 15562 -3772 15646 -3536
rect 15882 -3772 51326 -3536
rect 51562 -3772 51646 -3536
rect 51882 -3772 87326 -3536
rect 87562 -3772 87646 -3536
rect 87882 -3772 123326 -3536
rect 123562 -3772 123646 -3536
rect 123882 -3772 159326 -3536
rect 159562 -3772 159646 -3536
rect 159882 -3772 195326 -3536
rect 195562 -3772 195646 -3536
rect 195882 -3772 231326 -3536
rect 231562 -3772 231646 -3536
rect 231882 -3772 267326 -3536
rect 267562 -3772 267646 -3536
rect 267882 -3772 303326 -3536
rect 303562 -3772 303646 -3536
rect 303882 -3772 339326 -3536
rect 339562 -3772 339646 -3536
rect 339882 -3772 375326 -3536
rect 375562 -3772 375646 -3536
rect 375882 -3772 411326 -3536
rect 411562 -3772 411646 -3536
rect 411882 -3772 447326 -3536
rect 447562 -3772 447646 -3536
rect 447882 -3772 483326 -3536
rect 483562 -3772 483646 -3536
rect 483882 -3772 519326 -3536
rect 519562 -3772 519646 -3536
rect 519882 -3772 555326 -3536
rect 555562 -3772 555646 -3536
rect 555882 -3772 588532 -3536
rect 588768 -3772 588852 -3536
rect 589088 -3772 589120 -3536
rect -5196 -3856 589120 -3772
rect -5196 -4092 -5164 -3856
rect -4928 -4092 -4844 -3856
rect -4608 -4092 15326 -3856
rect 15562 -4092 15646 -3856
rect 15882 -4092 51326 -3856
rect 51562 -4092 51646 -3856
rect 51882 -4092 87326 -3856
rect 87562 -4092 87646 -3856
rect 87882 -4092 123326 -3856
rect 123562 -4092 123646 -3856
rect 123882 -4092 159326 -3856
rect 159562 -4092 159646 -3856
rect 159882 -4092 195326 -3856
rect 195562 -4092 195646 -3856
rect 195882 -4092 231326 -3856
rect 231562 -4092 231646 -3856
rect 231882 -4092 267326 -3856
rect 267562 -4092 267646 -3856
rect 267882 -4092 303326 -3856
rect 303562 -4092 303646 -3856
rect 303882 -4092 339326 -3856
rect 339562 -4092 339646 -3856
rect 339882 -4092 375326 -3856
rect 375562 -4092 375646 -3856
rect 375882 -4092 411326 -3856
rect 411562 -4092 411646 -3856
rect 411882 -4092 447326 -3856
rect 447562 -4092 447646 -3856
rect 447882 -4092 483326 -3856
rect 483562 -4092 483646 -3856
rect 483882 -4092 519326 -3856
rect 519562 -4092 519646 -3856
rect 519882 -4092 555326 -3856
rect 555562 -4092 555646 -3856
rect 555882 -4092 588532 -3856
rect 588768 -4092 588852 -3856
rect 589088 -4092 589120 -3856
rect -5196 -4124 589120 -4092
rect -6156 -4496 590080 -4464
rect -6156 -4732 -6124 -4496
rect -5888 -4732 -5804 -4496
rect -5568 -4732 19826 -4496
rect 20062 -4732 20146 -4496
rect 20382 -4732 55826 -4496
rect 56062 -4732 56146 -4496
rect 56382 -4732 91826 -4496
rect 92062 -4732 92146 -4496
rect 92382 -4732 127826 -4496
rect 128062 -4732 128146 -4496
rect 128382 -4732 163826 -4496
rect 164062 -4732 164146 -4496
rect 164382 -4732 199826 -4496
rect 200062 -4732 200146 -4496
rect 200382 -4732 235826 -4496
rect 236062 -4732 236146 -4496
rect 236382 -4732 271826 -4496
rect 272062 -4732 272146 -4496
rect 272382 -4732 307826 -4496
rect 308062 -4732 308146 -4496
rect 308382 -4732 343826 -4496
rect 344062 -4732 344146 -4496
rect 344382 -4732 379826 -4496
rect 380062 -4732 380146 -4496
rect 380382 -4732 415826 -4496
rect 416062 -4732 416146 -4496
rect 416382 -4732 451826 -4496
rect 452062 -4732 452146 -4496
rect 452382 -4732 487826 -4496
rect 488062 -4732 488146 -4496
rect 488382 -4732 523826 -4496
rect 524062 -4732 524146 -4496
rect 524382 -4732 559826 -4496
rect 560062 -4732 560146 -4496
rect 560382 -4732 589492 -4496
rect 589728 -4732 589812 -4496
rect 590048 -4732 590080 -4496
rect -6156 -4816 590080 -4732
rect -6156 -5052 -6124 -4816
rect -5888 -5052 -5804 -4816
rect -5568 -5052 19826 -4816
rect 20062 -5052 20146 -4816
rect 20382 -5052 55826 -4816
rect 56062 -5052 56146 -4816
rect 56382 -5052 91826 -4816
rect 92062 -5052 92146 -4816
rect 92382 -5052 127826 -4816
rect 128062 -5052 128146 -4816
rect 128382 -5052 163826 -4816
rect 164062 -5052 164146 -4816
rect 164382 -5052 199826 -4816
rect 200062 -5052 200146 -4816
rect 200382 -5052 235826 -4816
rect 236062 -5052 236146 -4816
rect 236382 -5052 271826 -4816
rect 272062 -5052 272146 -4816
rect 272382 -5052 307826 -4816
rect 308062 -5052 308146 -4816
rect 308382 -5052 343826 -4816
rect 344062 -5052 344146 -4816
rect 344382 -5052 379826 -4816
rect 380062 -5052 380146 -4816
rect 380382 -5052 415826 -4816
rect 416062 -5052 416146 -4816
rect 416382 -5052 451826 -4816
rect 452062 -5052 452146 -4816
rect 452382 -5052 487826 -4816
rect 488062 -5052 488146 -4816
rect 488382 -5052 523826 -4816
rect 524062 -5052 524146 -4816
rect 524382 -5052 559826 -4816
rect 560062 -5052 560146 -4816
rect 560382 -5052 589492 -4816
rect 589728 -5052 589812 -4816
rect 590048 -5052 590080 -4816
rect -6156 -5084 590080 -5052
rect -7116 -5456 591040 -5424
rect -7116 -5692 -7084 -5456
rect -6848 -5692 -6764 -5456
rect -6528 -5692 24326 -5456
rect 24562 -5692 24646 -5456
rect 24882 -5692 60326 -5456
rect 60562 -5692 60646 -5456
rect 60882 -5692 96326 -5456
rect 96562 -5692 96646 -5456
rect 96882 -5692 132326 -5456
rect 132562 -5692 132646 -5456
rect 132882 -5692 168326 -5456
rect 168562 -5692 168646 -5456
rect 168882 -5692 204326 -5456
rect 204562 -5692 204646 -5456
rect 204882 -5692 240326 -5456
rect 240562 -5692 240646 -5456
rect 240882 -5692 276326 -5456
rect 276562 -5692 276646 -5456
rect 276882 -5692 312326 -5456
rect 312562 -5692 312646 -5456
rect 312882 -5692 348326 -5456
rect 348562 -5692 348646 -5456
rect 348882 -5692 384326 -5456
rect 384562 -5692 384646 -5456
rect 384882 -5692 420326 -5456
rect 420562 -5692 420646 -5456
rect 420882 -5692 456326 -5456
rect 456562 -5692 456646 -5456
rect 456882 -5692 492326 -5456
rect 492562 -5692 492646 -5456
rect 492882 -5692 528326 -5456
rect 528562 -5692 528646 -5456
rect 528882 -5692 564326 -5456
rect 564562 -5692 564646 -5456
rect 564882 -5692 590452 -5456
rect 590688 -5692 590772 -5456
rect 591008 -5692 591040 -5456
rect -7116 -5776 591040 -5692
rect -7116 -6012 -7084 -5776
rect -6848 -6012 -6764 -5776
rect -6528 -6012 24326 -5776
rect 24562 -6012 24646 -5776
rect 24882 -6012 60326 -5776
rect 60562 -6012 60646 -5776
rect 60882 -6012 96326 -5776
rect 96562 -6012 96646 -5776
rect 96882 -6012 132326 -5776
rect 132562 -6012 132646 -5776
rect 132882 -6012 168326 -5776
rect 168562 -6012 168646 -5776
rect 168882 -6012 204326 -5776
rect 204562 -6012 204646 -5776
rect 204882 -6012 240326 -5776
rect 240562 -6012 240646 -5776
rect 240882 -6012 276326 -5776
rect 276562 -6012 276646 -5776
rect 276882 -6012 312326 -5776
rect 312562 -6012 312646 -5776
rect 312882 -6012 348326 -5776
rect 348562 -6012 348646 -5776
rect 348882 -6012 384326 -5776
rect 384562 -6012 384646 -5776
rect 384882 -6012 420326 -5776
rect 420562 -6012 420646 -5776
rect 420882 -6012 456326 -5776
rect 456562 -6012 456646 -5776
rect 456882 -6012 492326 -5776
rect 492562 -6012 492646 -5776
rect 492882 -6012 528326 -5776
rect 528562 -6012 528646 -5776
rect 528882 -6012 564326 -5776
rect 564562 -6012 564646 -5776
rect 564882 -6012 590452 -5776
rect 590688 -6012 590772 -5776
rect 591008 -6012 591040 -5776
rect -7116 -6044 591040 -6012
rect -8076 -6416 592000 -6384
rect -8076 -6652 -8044 -6416
rect -7808 -6652 -7724 -6416
rect -7488 -6652 28826 -6416
rect 29062 -6652 29146 -6416
rect 29382 -6652 64826 -6416
rect 65062 -6652 65146 -6416
rect 65382 -6652 100826 -6416
rect 101062 -6652 101146 -6416
rect 101382 -6652 136826 -6416
rect 137062 -6652 137146 -6416
rect 137382 -6652 172826 -6416
rect 173062 -6652 173146 -6416
rect 173382 -6652 208826 -6416
rect 209062 -6652 209146 -6416
rect 209382 -6652 244826 -6416
rect 245062 -6652 245146 -6416
rect 245382 -6652 280826 -6416
rect 281062 -6652 281146 -6416
rect 281382 -6652 316826 -6416
rect 317062 -6652 317146 -6416
rect 317382 -6652 352826 -6416
rect 353062 -6652 353146 -6416
rect 353382 -6652 388826 -6416
rect 389062 -6652 389146 -6416
rect 389382 -6652 424826 -6416
rect 425062 -6652 425146 -6416
rect 425382 -6652 460826 -6416
rect 461062 -6652 461146 -6416
rect 461382 -6652 496826 -6416
rect 497062 -6652 497146 -6416
rect 497382 -6652 532826 -6416
rect 533062 -6652 533146 -6416
rect 533382 -6652 568826 -6416
rect 569062 -6652 569146 -6416
rect 569382 -6652 591412 -6416
rect 591648 -6652 591732 -6416
rect 591968 -6652 592000 -6416
rect -8076 -6736 592000 -6652
rect -8076 -6972 -8044 -6736
rect -7808 -6972 -7724 -6736
rect -7488 -6972 28826 -6736
rect 29062 -6972 29146 -6736
rect 29382 -6972 64826 -6736
rect 65062 -6972 65146 -6736
rect 65382 -6972 100826 -6736
rect 101062 -6972 101146 -6736
rect 101382 -6972 136826 -6736
rect 137062 -6972 137146 -6736
rect 137382 -6972 172826 -6736
rect 173062 -6972 173146 -6736
rect 173382 -6972 208826 -6736
rect 209062 -6972 209146 -6736
rect 209382 -6972 244826 -6736
rect 245062 -6972 245146 -6736
rect 245382 -6972 280826 -6736
rect 281062 -6972 281146 -6736
rect 281382 -6972 316826 -6736
rect 317062 -6972 317146 -6736
rect 317382 -6972 352826 -6736
rect 353062 -6972 353146 -6736
rect 353382 -6972 388826 -6736
rect 389062 -6972 389146 -6736
rect 389382 -6972 424826 -6736
rect 425062 -6972 425146 -6736
rect 425382 -6972 460826 -6736
rect 461062 -6972 461146 -6736
rect 461382 -6972 496826 -6736
rect 497062 -6972 497146 -6736
rect 497382 -6972 532826 -6736
rect 533062 -6972 533146 -6736
rect 533382 -6972 568826 -6736
rect 569062 -6972 569146 -6736
rect 569382 -6972 591412 -6736
rect 591648 -6972 591732 -6736
rect 591968 -6972 592000 -6736
rect -8076 -7004 592000 -6972
rect -9036 -7376 592960 -7344
rect -9036 -7612 -9004 -7376
rect -8768 -7612 -8684 -7376
rect -8448 -7612 33326 -7376
rect 33562 -7612 33646 -7376
rect 33882 -7612 69326 -7376
rect 69562 -7612 69646 -7376
rect 69882 -7612 105326 -7376
rect 105562 -7612 105646 -7376
rect 105882 -7612 141326 -7376
rect 141562 -7612 141646 -7376
rect 141882 -7612 177326 -7376
rect 177562 -7612 177646 -7376
rect 177882 -7612 213326 -7376
rect 213562 -7612 213646 -7376
rect 213882 -7612 249326 -7376
rect 249562 -7612 249646 -7376
rect 249882 -7612 285326 -7376
rect 285562 -7612 285646 -7376
rect 285882 -7612 321326 -7376
rect 321562 -7612 321646 -7376
rect 321882 -7612 357326 -7376
rect 357562 -7612 357646 -7376
rect 357882 -7612 393326 -7376
rect 393562 -7612 393646 -7376
rect 393882 -7612 429326 -7376
rect 429562 -7612 429646 -7376
rect 429882 -7612 465326 -7376
rect 465562 -7612 465646 -7376
rect 465882 -7612 501326 -7376
rect 501562 -7612 501646 -7376
rect 501882 -7612 537326 -7376
rect 537562 -7612 537646 -7376
rect 537882 -7612 573326 -7376
rect 573562 -7612 573646 -7376
rect 573882 -7612 592372 -7376
rect 592608 -7612 592692 -7376
rect 592928 -7612 592960 -7376
rect -9036 -7696 592960 -7612
rect -9036 -7932 -9004 -7696
rect -8768 -7932 -8684 -7696
rect -8448 -7932 33326 -7696
rect 33562 -7932 33646 -7696
rect 33882 -7932 69326 -7696
rect 69562 -7932 69646 -7696
rect 69882 -7932 105326 -7696
rect 105562 -7932 105646 -7696
rect 105882 -7932 141326 -7696
rect 141562 -7932 141646 -7696
rect 141882 -7932 177326 -7696
rect 177562 -7932 177646 -7696
rect 177882 -7932 213326 -7696
rect 213562 -7932 213646 -7696
rect 213882 -7932 249326 -7696
rect 249562 -7932 249646 -7696
rect 249882 -7932 285326 -7696
rect 285562 -7932 285646 -7696
rect 285882 -7932 321326 -7696
rect 321562 -7932 321646 -7696
rect 321882 -7932 357326 -7696
rect 357562 -7932 357646 -7696
rect 357882 -7932 393326 -7696
rect 393562 -7932 393646 -7696
rect 393882 -7932 429326 -7696
rect 429562 -7932 429646 -7696
rect 429882 -7932 465326 -7696
rect 465562 -7932 465646 -7696
rect 465882 -7932 501326 -7696
rect 501562 -7932 501646 -7696
rect 501882 -7932 537326 -7696
rect 537562 -7932 537646 -7696
rect 537882 -7932 573326 -7696
rect 573562 -7932 573646 -7696
rect 573882 -7932 592372 -7696
rect 592608 -7932 592692 -7696
rect 592928 -7932 592960 -7696
rect -9036 -7964 592960 -7932
use macro_7  u_macro_7
timestamp 0
transform 1 0 80000 0 1 100000
box 1066 0 48890 50000
<< labels >>
flabel metal3 s 583520 7700 584960 7940 0 FreeSans 960 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 583520 476900 584960 477140 0 FreeSans 960 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 583520 523820 584960 524060 0 FreeSans 960 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 583520 570740 584960 570980 0 FreeSans 960 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 583520 617660 584960 617900 0 FreeSans 960 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 583520 664580 584960 664820 0 FreeSans 960 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 572966 703520 573078 704960 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 508106 703520 508218 704960 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 443246 703520 443358 704960 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 378386 703520 378498 704960 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 313526 703520 313638 704960 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 583520 54620 584960 54860 0 FreeSans 960 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 248666 703520 248778 704960 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 183806 703520 183918 704960 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 118946 703520 119058 704960 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 54086 703520 54198 704960 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 694772 480 695012 0 FreeSans 960 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 644588 480 644828 0 FreeSans 960 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 594404 480 594644 0 FreeSans 960 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 544220 480 544460 0 FreeSans 960 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 494036 480 494276 0 FreeSans 960 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 443852 480 444092 0 FreeSans 960 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 583520 101540 584960 101780 0 FreeSans 960 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 393668 480 393908 0 FreeSans 960 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 343484 480 343724 0 FreeSans 960 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 293300 480 293540 0 FreeSans 960 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 243116 480 243356 0 FreeSans 960 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 192932 480 193172 0 FreeSans 960 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 142748 480 142988 0 FreeSans 960 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 92564 480 92804 0 FreeSans 960 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 42380 480 42620 0 FreeSans 960 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 583520 148460 584960 148700 0 FreeSans 960 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 583520 195380 584960 195620 0 FreeSans 960 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 583520 242300 584960 242540 0 FreeSans 960 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 583520 289220 584960 289460 0 FreeSans 960 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 583520 336140 584960 336380 0 FreeSans 960 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 583520 383060 584960 383300 0 FreeSans 960 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 583520 429980 584960 430220 0 FreeSans 960 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 583520 38980 584960 39220 0 FreeSans 960 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 583520 508180 584960 508420 0 FreeSans 960 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 583520 555100 584960 555340 0 FreeSans 960 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 583520 602020 584960 602260 0 FreeSans 960 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 583520 648940 584960 649180 0 FreeSans 960 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 583520 695860 584960 696100 0 FreeSans 960 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 529726 703520 529838 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 464866 703520 464978 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 400006 703520 400118 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 335146 703520 335258 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 270286 703520 270398 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 583520 85900 584960 86140 0 FreeSans 960 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 205426 703520 205538 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 140566 703520 140678 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 75706 703520 75818 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 10846 703520 10958 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 661316 480 661556 0 FreeSans 960 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 611132 480 611372 0 FreeSans 960 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 560948 480 561188 0 FreeSans 960 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 510764 480 511004 0 FreeSans 960 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 460580 480 460820 0 FreeSans 960 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 583520 132820 584960 133060 0 FreeSans 960 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 360212 480 360452 0 FreeSans 960 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 310028 480 310268 0 FreeSans 960 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 259844 480 260084 0 FreeSans 960 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 209660 480 209900 0 FreeSans 960 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 159476 480 159716 0 FreeSans 960 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 109292 480 109532 0 FreeSans 960 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 59108 480 59348 0 FreeSans 960 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8924 480 9164 0 FreeSans 960 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 583520 179740 584960 179980 0 FreeSans 960 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 583520 226660 584960 226900 0 FreeSans 960 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 583520 273580 584960 273820 0 FreeSans 960 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 583520 320500 584960 320740 0 FreeSans 960 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 583520 367420 584960 367660 0 FreeSans 960 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 583520 414340 584960 414580 0 FreeSans 960 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 583520 461260 584960 461500 0 FreeSans 960 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 583520 23340 584960 23580 0 FreeSans 960 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 583520 492540 584960 492780 0 FreeSans 960 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 583520 539460 584960 539700 0 FreeSans 960 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 583520 586380 584960 586620 0 FreeSans 960 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 583520 633300 584960 633540 0 FreeSans 960 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 583520 680220 584960 680460 0 FreeSans 960 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 551346 703520 551458 704960 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 486486 703520 486598 704960 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 421626 703520 421738 704960 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 356766 703520 356878 704960 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 291906 703520 292018 704960 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 583520 70260 584960 70500 0 FreeSans 960 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 227046 703520 227158 704960 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 162186 703520 162298 704960 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 97326 703520 97438 704960 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 32466 703520 32578 704960 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 678044 480 678284 0 FreeSans 960 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 627860 480 628100 0 FreeSans 960 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 577676 480 577916 0 FreeSans 960 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 527492 480 527732 0 FreeSans 960 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 477308 480 477548 0 FreeSans 960 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 427124 480 427364 0 FreeSans 960 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 583520 117180 584960 117420 0 FreeSans 960 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 376940 480 377180 0 FreeSans 960 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 326756 480 326996 0 FreeSans 960 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 276572 480 276812 0 FreeSans 960 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 226388 480 226628 0 FreeSans 960 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 176204 480 176444 0 FreeSans 960 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 126020 480 126260 0 FreeSans 960 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 75836 480 76076 0 FreeSans 960 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 25652 480 25892 0 FreeSans 960 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 583520 164100 584960 164340 0 FreeSans 960 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 583520 211020 584960 211260 0 FreeSans 960 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 583520 257940 584960 258180 0 FreeSans 960 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 583520 304860 584960 305100 0 FreeSans 960 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 583520 398700 584960 398940 0 FreeSans 960 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 583520 445620 584960 445860 0 FreeSans 960 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 139002 -960 139114 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 470202 -960 470314 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 115 nsew signal input
flabel metal2 s 473514 -960 473626 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 116 nsew signal input
flabel metal2 s 476826 -960 476938 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 117 nsew signal input
flabel metal2 s 480138 -960 480250 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 118 nsew signal input
flabel metal2 s 483450 -960 483562 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 119 nsew signal input
flabel metal2 s 486762 -960 486874 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 120 nsew signal input
flabel metal2 s 490074 -960 490186 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 121 nsew signal input
flabel metal2 s 493386 -960 493498 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 122 nsew signal input
flabel metal2 s 496698 -960 496810 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 123 nsew signal input
flabel metal2 s 500010 -960 500122 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 124 nsew signal input
flabel metal2 s 172122 -960 172234 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 125 nsew signal input
flabel metal2 s 503322 -960 503434 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 126 nsew signal input
flabel metal2 s 506634 -960 506746 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 127 nsew signal input
flabel metal2 s 509946 -960 510058 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 128 nsew signal input
flabel metal2 s 513258 -960 513370 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 129 nsew signal input
flabel metal2 s 516570 -960 516682 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 130 nsew signal input
flabel metal2 s 519882 -960 519994 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 131 nsew signal input
flabel metal2 s 523194 -960 523306 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 132 nsew signal input
flabel metal2 s 526506 -960 526618 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 133 nsew signal input
flabel metal2 s 529818 -960 529930 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 134 nsew signal input
flabel metal2 s 533130 -960 533242 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 135 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 136 nsew signal input
flabel metal2 s 536442 -960 536554 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 137 nsew signal input
flabel metal2 s 539754 -960 539866 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 138 nsew signal input
flabel metal2 s 543066 -960 543178 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 139 nsew signal input
flabel metal2 s 546378 -960 546490 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 140 nsew signal input
flabel metal2 s 549690 -960 549802 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 141 nsew signal input
flabel metal2 s 553002 -960 553114 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 142 nsew signal input
flabel metal2 s 556314 -960 556426 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 143 nsew signal input
flabel metal2 s 559626 -960 559738 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 144 nsew signal input
flabel metal2 s 178746 -960 178858 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 145 nsew signal input
flabel metal2 s 182058 -960 182170 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 146 nsew signal input
flabel metal2 s 185370 -960 185482 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 147 nsew signal input
flabel metal2 s 188682 -960 188794 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 148 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 149 nsew signal input
flabel metal2 s 195306 -960 195418 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 150 nsew signal input
flabel metal2 s 198618 -960 198730 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 151 nsew signal input
flabel metal2 s 201930 -960 202042 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 152 nsew signal input
flabel metal2 s 142314 -960 142426 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 153 nsew signal input
flabel metal2 s 205242 -960 205354 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 154 nsew signal input
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 155 nsew signal input
flabel metal2 s 211866 -960 211978 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 156 nsew signal input
flabel metal2 s 215178 -960 215290 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 157 nsew signal input
flabel metal2 s 218490 -960 218602 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 158 nsew signal input
flabel metal2 s 221802 -960 221914 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 159 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 160 nsew signal input
flabel metal2 s 228426 -960 228538 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 161 nsew signal input
flabel metal2 s 231738 -960 231850 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 162 nsew signal input
flabel metal2 s 235050 -960 235162 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 163 nsew signal input
flabel metal2 s 145626 -960 145738 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 164 nsew signal input
flabel metal2 s 238362 -960 238474 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 165 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 166 nsew signal input
flabel metal2 s 244986 -960 245098 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 167 nsew signal input
flabel metal2 s 248298 -960 248410 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 168 nsew signal input
flabel metal2 s 251610 -960 251722 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 169 nsew signal input
flabel metal2 s 254922 -960 255034 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 170 nsew signal input
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 171 nsew signal input
flabel metal2 s 261546 -960 261658 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 172 nsew signal input
flabel metal2 s 264858 -960 264970 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 173 nsew signal input
flabel metal2 s 268170 -960 268282 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 174 nsew signal input
flabel metal2 s 148938 -960 149050 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 175 nsew signal input
flabel metal2 s 271482 -960 271594 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 176 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 177 nsew signal input
flabel metal2 s 278106 -960 278218 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 178 nsew signal input
flabel metal2 s 281418 -960 281530 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 179 nsew signal input
flabel metal2 s 284730 -960 284842 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 180 nsew signal input
flabel metal2 s 288042 -960 288154 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 181 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 182 nsew signal input
flabel metal2 s 294666 -960 294778 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 183 nsew signal input
flabel metal2 s 297978 -960 298090 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 184 nsew signal input
flabel metal2 s 301290 -960 301402 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 185 nsew signal input
flabel metal2 s 152250 -960 152362 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 186 nsew signal input
flabel metal2 s 304602 -960 304714 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 187 nsew signal input
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 188 nsew signal input
flabel metal2 s 311226 -960 311338 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 189 nsew signal input
flabel metal2 s 314538 -960 314650 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 190 nsew signal input
flabel metal2 s 317850 -960 317962 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 191 nsew signal input
flabel metal2 s 321162 -960 321274 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 192 nsew signal input
flabel metal2 s 324474 -960 324586 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 193 nsew signal input
flabel metal2 s 327786 -960 327898 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 194 nsew signal input
flabel metal2 s 331098 -960 331210 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 195 nsew signal input
flabel metal2 s 334410 -960 334522 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 196 nsew signal input
flabel metal2 s 155562 -960 155674 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 197 nsew signal input
flabel metal2 s 337722 -960 337834 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 198 nsew signal input
flabel metal2 s 341034 -960 341146 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 199 nsew signal input
flabel metal2 s 344346 -960 344458 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 200 nsew signal input
flabel metal2 s 347658 -960 347770 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 201 nsew signal input
flabel metal2 s 350970 -960 351082 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 202 nsew signal input
flabel metal2 s 354282 -960 354394 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 203 nsew signal input
flabel metal2 s 357594 -960 357706 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 204 nsew signal input
flabel metal2 s 360906 -960 361018 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 205 nsew signal input
flabel metal2 s 364218 -960 364330 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 206 nsew signal input
flabel metal2 s 367530 -960 367642 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 207 nsew signal input
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 208 nsew signal input
flabel metal2 s 370842 -960 370954 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 209 nsew signal input
flabel metal2 s 374154 -960 374266 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 210 nsew signal input
flabel metal2 s 377466 -960 377578 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 211 nsew signal input
flabel metal2 s 380778 -960 380890 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 212 nsew signal input
flabel metal2 s 384090 -960 384202 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 213 nsew signal input
flabel metal2 s 387402 -960 387514 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 214 nsew signal input
flabel metal2 s 390714 -960 390826 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 215 nsew signal input
flabel metal2 s 394026 -960 394138 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 216 nsew signal input
flabel metal2 s 397338 -960 397450 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 217 nsew signal input
flabel metal2 s 400650 -960 400762 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 218 nsew signal input
flabel metal2 s 162186 -960 162298 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 219 nsew signal input
flabel metal2 s 403962 -960 404074 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 220 nsew signal input
flabel metal2 s 407274 -960 407386 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 221 nsew signal input
flabel metal2 s 410586 -960 410698 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 222 nsew signal input
flabel metal2 s 413898 -960 414010 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 223 nsew signal input
flabel metal2 s 417210 -960 417322 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 224 nsew signal input
flabel metal2 s 420522 -960 420634 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 225 nsew signal input
flabel metal2 s 423834 -960 423946 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 226 nsew signal input
flabel metal2 s 427146 -960 427258 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 227 nsew signal input
flabel metal2 s 430458 -960 430570 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 228 nsew signal input
flabel metal2 s 433770 -960 433882 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 229 nsew signal input
flabel metal2 s 165498 -960 165610 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 230 nsew signal input
flabel metal2 s 437082 -960 437194 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 231 nsew signal input
flabel metal2 s 440394 -960 440506 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 232 nsew signal input
flabel metal2 s 443706 -960 443818 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 233 nsew signal input
flabel metal2 s 447018 -960 447130 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 234 nsew signal input
flabel metal2 s 450330 -960 450442 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 235 nsew signal input
flabel metal2 s 453642 -960 453754 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 236 nsew signal input
flabel metal2 s 456954 -960 457066 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 237 nsew signal input
flabel metal2 s 460266 -960 460378 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 238 nsew signal input
flabel metal2 s 463578 -960 463690 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 239 nsew signal input
flabel metal2 s 466890 -960 467002 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 240 nsew signal input
flabel metal2 s 168810 -960 168922 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 241 nsew signal input
flabel metal2 s 140106 -960 140218 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 242 nsew signal tristate
flabel metal2 s 471306 -960 471418 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 243 nsew signal tristate
flabel metal2 s 474618 -960 474730 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 244 nsew signal tristate
flabel metal2 s 477930 -960 478042 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 245 nsew signal tristate
flabel metal2 s 481242 -960 481354 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 246 nsew signal tristate
flabel metal2 s 484554 -960 484666 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 247 nsew signal tristate
flabel metal2 s 487866 -960 487978 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 248 nsew signal tristate
flabel metal2 s 491178 -960 491290 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 249 nsew signal tristate
flabel metal2 s 494490 -960 494602 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 250 nsew signal tristate
flabel metal2 s 497802 -960 497914 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 251 nsew signal tristate
flabel metal2 s 501114 -960 501226 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 252 nsew signal tristate
flabel metal2 s 173226 -960 173338 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 253 nsew signal tristate
flabel metal2 s 504426 -960 504538 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 254 nsew signal tristate
flabel metal2 s 507738 -960 507850 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 255 nsew signal tristate
flabel metal2 s 511050 -960 511162 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 256 nsew signal tristate
flabel metal2 s 514362 -960 514474 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 257 nsew signal tristate
flabel metal2 s 517674 -960 517786 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 258 nsew signal tristate
flabel metal2 s 520986 -960 521098 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 259 nsew signal tristate
flabel metal2 s 524298 -960 524410 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 260 nsew signal tristate
flabel metal2 s 527610 -960 527722 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 261 nsew signal tristate
flabel metal2 s 530922 -960 531034 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 262 nsew signal tristate
flabel metal2 s 534234 -960 534346 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 263 nsew signal tristate
flabel metal2 s 176538 -960 176650 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 264 nsew signal tristate
flabel metal2 s 537546 -960 537658 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 265 nsew signal tristate
flabel metal2 s 540858 -960 540970 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 266 nsew signal tristate
flabel metal2 s 544170 -960 544282 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 267 nsew signal tristate
flabel metal2 s 547482 -960 547594 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 268 nsew signal tristate
flabel metal2 s 550794 -960 550906 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 269 nsew signal tristate
flabel metal2 s 554106 -960 554218 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 270 nsew signal tristate
flabel metal2 s 557418 -960 557530 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 271 nsew signal tristate
flabel metal2 s 560730 -960 560842 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 272 nsew signal tristate
flabel metal2 s 179850 -960 179962 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 273 nsew signal tristate
flabel metal2 s 183162 -960 183274 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 274 nsew signal tristate
flabel metal2 s 186474 -960 186586 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 275 nsew signal tristate
flabel metal2 s 189786 -960 189898 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 276 nsew signal tristate
flabel metal2 s 193098 -960 193210 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 277 nsew signal tristate
flabel metal2 s 196410 -960 196522 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 278 nsew signal tristate
flabel metal2 s 199722 -960 199834 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 279 nsew signal tristate
flabel metal2 s 203034 -960 203146 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 280 nsew signal tristate
flabel metal2 s 143418 -960 143530 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 281 nsew signal tristate
flabel metal2 s 206346 -960 206458 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 282 nsew signal tristate
flabel metal2 s 209658 -960 209770 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 283 nsew signal tristate
flabel metal2 s 212970 -960 213082 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 284 nsew signal tristate
flabel metal2 s 216282 -960 216394 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 285 nsew signal tristate
flabel metal2 s 219594 -960 219706 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 286 nsew signal tristate
flabel metal2 s 222906 -960 223018 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 287 nsew signal tristate
flabel metal2 s 226218 -960 226330 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 288 nsew signal tristate
flabel metal2 s 229530 -960 229642 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 289 nsew signal tristate
flabel metal2 s 232842 -960 232954 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 290 nsew signal tristate
flabel metal2 s 236154 -960 236266 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 291 nsew signal tristate
flabel metal2 s 146730 -960 146842 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 292 nsew signal tristate
flabel metal2 s 239466 -960 239578 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 293 nsew signal tristate
flabel metal2 s 242778 -960 242890 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 294 nsew signal tristate
flabel metal2 s 246090 -960 246202 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 295 nsew signal tristate
flabel metal2 s 249402 -960 249514 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 296 nsew signal tristate
flabel metal2 s 252714 -960 252826 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 297 nsew signal tristate
flabel metal2 s 256026 -960 256138 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 298 nsew signal tristate
flabel metal2 s 259338 -960 259450 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 299 nsew signal tristate
flabel metal2 s 262650 -960 262762 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 300 nsew signal tristate
flabel metal2 s 265962 -960 266074 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 301 nsew signal tristate
flabel metal2 s 269274 -960 269386 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 302 nsew signal tristate
flabel metal2 s 150042 -960 150154 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 303 nsew signal tristate
flabel metal2 s 272586 -960 272698 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 304 nsew signal tristate
flabel metal2 s 275898 -960 276010 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 305 nsew signal tristate
flabel metal2 s 279210 -960 279322 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 306 nsew signal tristate
flabel metal2 s 282522 -960 282634 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 307 nsew signal tristate
flabel metal2 s 285834 -960 285946 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 308 nsew signal tristate
flabel metal2 s 289146 -960 289258 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 309 nsew signal tristate
flabel metal2 s 292458 -960 292570 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 310 nsew signal tristate
flabel metal2 s 295770 -960 295882 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 311 nsew signal tristate
flabel metal2 s 299082 -960 299194 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 312 nsew signal tristate
flabel metal2 s 302394 -960 302506 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 313 nsew signal tristate
flabel metal2 s 153354 -960 153466 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 314 nsew signal tristate
flabel metal2 s 305706 -960 305818 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 315 nsew signal tristate
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 316 nsew signal tristate
flabel metal2 s 312330 -960 312442 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 317 nsew signal tristate
flabel metal2 s 315642 -960 315754 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 318 nsew signal tristate
flabel metal2 s 318954 -960 319066 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 319 nsew signal tristate
flabel metal2 s 322266 -960 322378 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 320 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 321 nsew signal tristate
flabel metal2 s 328890 -960 329002 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 322 nsew signal tristate
flabel metal2 s 332202 -960 332314 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 323 nsew signal tristate
flabel metal2 s 335514 -960 335626 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 324 nsew signal tristate
flabel metal2 s 156666 -960 156778 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 325 nsew signal tristate
flabel metal2 s 338826 -960 338938 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 326 nsew signal tristate
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 327 nsew signal tristate
flabel metal2 s 345450 -960 345562 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 328 nsew signal tristate
flabel metal2 s 348762 -960 348874 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 329 nsew signal tristate
flabel metal2 s 352074 -960 352186 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 330 nsew signal tristate
flabel metal2 s 355386 -960 355498 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 331 nsew signal tristate
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 332 nsew signal tristate
flabel metal2 s 362010 -960 362122 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 333 nsew signal tristate
flabel metal2 s 365322 -960 365434 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 334 nsew signal tristate
flabel metal2 s 368634 -960 368746 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 335 nsew signal tristate
flabel metal2 s 159978 -960 160090 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 336 nsew signal tristate
flabel metal2 s 371946 -960 372058 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 337 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 338 nsew signal tristate
flabel metal2 s 378570 -960 378682 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 339 nsew signal tristate
flabel metal2 s 381882 -960 381994 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 340 nsew signal tristate
flabel metal2 s 385194 -960 385306 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 341 nsew signal tristate
flabel metal2 s 388506 -960 388618 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 342 nsew signal tristate
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 343 nsew signal tristate
flabel metal2 s 395130 -960 395242 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 344 nsew signal tristate
flabel metal2 s 398442 -960 398554 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 345 nsew signal tristate
flabel metal2 s 401754 -960 401866 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 346 nsew signal tristate
flabel metal2 s 163290 -960 163402 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 347 nsew signal tristate
flabel metal2 s 405066 -960 405178 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 348 nsew signal tristate
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 349 nsew signal tristate
flabel metal2 s 411690 -960 411802 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 350 nsew signal tristate
flabel metal2 s 415002 -960 415114 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 351 nsew signal tristate
flabel metal2 s 418314 -960 418426 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 352 nsew signal tristate
flabel metal2 s 421626 -960 421738 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 353 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 354 nsew signal tristate
flabel metal2 s 428250 -960 428362 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 355 nsew signal tristate
flabel metal2 s 431562 -960 431674 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 356 nsew signal tristate
flabel metal2 s 434874 -960 434986 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 357 nsew signal tristate
flabel metal2 s 166602 -960 166714 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 358 nsew signal tristate
flabel metal2 s 438186 -960 438298 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 359 nsew signal tristate
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 360 nsew signal tristate
flabel metal2 s 444810 -960 444922 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 361 nsew signal tristate
flabel metal2 s 448122 -960 448234 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 362 nsew signal tristate
flabel metal2 s 451434 -960 451546 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 363 nsew signal tristate
flabel metal2 s 454746 -960 454858 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 364 nsew signal tristate
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 365 nsew signal tristate
flabel metal2 s 461370 -960 461482 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 366 nsew signal tristate
flabel metal2 s 464682 -960 464794 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 367 nsew signal tristate
flabel metal2 s 467994 -960 468106 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 368 nsew signal tristate
flabel metal2 s 169914 -960 170026 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 369 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 370 nsew signal input
flabel metal2 s 472410 -960 472522 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 371 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 372 nsew signal input
flabel metal2 s 479034 -960 479146 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 373 nsew signal input
flabel metal2 s 482346 -960 482458 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 374 nsew signal input
flabel metal2 s 485658 -960 485770 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 375 nsew signal input
flabel metal2 s 488970 -960 489082 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 376 nsew signal input
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 377 nsew signal input
flabel metal2 s 495594 -960 495706 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 378 nsew signal input
flabel metal2 s 498906 -960 499018 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 379 nsew signal input
flabel metal2 s 502218 -960 502330 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 380 nsew signal input
flabel metal2 s 174330 -960 174442 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 381 nsew signal input
flabel metal2 s 505530 -960 505642 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 382 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 383 nsew signal input
flabel metal2 s 512154 -960 512266 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 384 nsew signal input
flabel metal2 s 515466 -960 515578 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 385 nsew signal input
flabel metal2 s 518778 -960 518890 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 386 nsew signal input
flabel metal2 s 522090 -960 522202 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 387 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 388 nsew signal input
flabel metal2 s 528714 -960 528826 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 389 nsew signal input
flabel metal2 s 532026 -960 532138 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 390 nsew signal input
flabel metal2 s 535338 -960 535450 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 391 nsew signal input
flabel metal2 s 177642 -960 177754 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 392 nsew signal input
flabel metal2 s 538650 -960 538762 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 393 nsew signal input
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 394 nsew signal input
flabel metal2 s 545274 -960 545386 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 395 nsew signal input
flabel metal2 s 548586 -960 548698 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 396 nsew signal input
flabel metal2 s 551898 -960 552010 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 397 nsew signal input
flabel metal2 s 555210 -960 555322 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 398 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 399 nsew signal input
flabel metal2 s 561834 -960 561946 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 400 nsew signal input
flabel metal2 s 180954 -960 181066 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 401 nsew signal input
flabel metal2 s 184266 -960 184378 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 402 nsew signal input
flabel metal2 s 187578 -960 187690 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 403 nsew signal input
flabel metal2 s 190890 -960 191002 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 404 nsew signal input
flabel metal2 s 194202 -960 194314 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 405 nsew signal input
flabel metal2 s 197514 -960 197626 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 406 nsew signal input
flabel metal2 s 200826 -960 200938 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 407 nsew signal input
flabel metal2 s 204138 -960 204250 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 408 nsew signal input
flabel metal2 s 144522 -960 144634 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 409 nsew signal input
flabel metal2 s 207450 -960 207562 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 410 nsew signal input
flabel metal2 s 210762 -960 210874 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 411 nsew signal input
flabel metal2 s 214074 -960 214186 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 412 nsew signal input
flabel metal2 s 217386 -960 217498 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 413 nsew signal input
flabel metal2 s 220698 -960 220810 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 414 nsew signal input
flabel metal2 s 224010 -960 224122 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 415 nsew signal input
flabel metal2 s 227322 -960 227434 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 416 nsew signal input
flabel metal2 s 230634 -960 230746 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 417 nsew signal input
flabel metal2 s 233946 -960 234058 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 418 nsew signal input
flabel metal2 s 237258 -960 237370 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 419 nsew signal input
flabel metal2 s 147834 -960 147946 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 420 nsew signal input
flabel metal2 s 240570 -960 240682 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 421 nsew signal input
flabel metal2 s 243882 -960 243994 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 422 nsew signal input
flabel metal2 s 247194 -960 247306 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 423 nsew signal input
flabel metal2 s 250506 -960 250618 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 424 nsew signal input
flabel metal2 s 253818 -960 253930 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 425 nsew signal input
flabel metal2 s 257130 -960 257242 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 426 nsew signal input
flabel metal2 s 260442 -960 260554 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 427 nsew signal input
flabel metal2 s 263754 -960 263866 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 428 nsew signal input
flabel metal2 s 267066 -960 267178 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 429 nsew signal input
flabel metal2 s 270378 -960 270490 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 430 nsew signal input
flabel metal2 s 151146 -960 151258 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 431 nsew signal input
flabel metal2 s 273690 -960 273802 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 432 nsew signal input
flabel metal2 s 277002 -960 277114 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 433 nsew signal input
flabel metal2 s 280314 -960 280426 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 434 nsew signal input
flabel metal2 s 283626 -960 283738 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 435 nsew signal input
flabel metal2 s 286938 -960 287050 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 436 nsew signal input
flabel metal2 s 290250 -960 290362 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 437 nsew signal input
flabel metal2 s 293562 -960 293674 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 438 nsew signal input
flabel metal2 s 296874 -960 296986 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 439 nsew signal input
flabel metal2 s 300186 -960 300298 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 440 nsew signal input
flabel metal2 s 303498 -960 303610 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 441 nsew signal input
flabel metal2 s 154458 -960 154570 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 442 nsew signal input
flabel metal2 s 306810 -960 306922 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 443 nsew signal input
flabel metal2 s 310122 -960 310234 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 444 nsew signal input
flabel metal2 s 313434 -960 313546 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 445 nsew signal input
flabel metal2 s 316746 -960 316858 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 446 nsew signal input
flabel metal2 s 320058 -960 320170 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 447 nsew signal input
flabel metal2 s 323370 -960 323482 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 448 nsew signal input
flabel metal2 s 326682 -960 326794 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 449 nsew signal input
flabel metal2 s 329994 -960 330106 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 450 nsew signal input
flabel metal2 s 333306 -960 333418 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 451 nsew signal input
flabel metal2 s 336618 -960 336730 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 452 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 453 nsew signal input
flabel metal2 s 339930 -960 340042 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 454 nsew signal input
flabel metal2 s 343242 -960 343354 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 455 nsew signal input
flabel metal2 s 346554 -960 346666 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 456 nsew signal input
flabel metal2 s 349866 -960 349978 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 457 nsew signal input
flabel metal2 s 353178 -960 353290 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 458 nsew signal input
flabel metal2 s 356490 -960 356602 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 459 nsew signal input
flabel metal2 s 359802 -960 359914 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 460 nsew signal input
flabel metal2 s 363114 -960 363226 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 461 nsew signal input
flabel metal2 s 366426 -960 366538 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 462 nsew signal input
flabel metal2 s 369738 -960 369850 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 463 nsew signal input
flabel metal2 s 161082 -960 161194 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 464 nsew signal input
flabel metal2 s 373050 -960 373162 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 465 nsew signal input
flabel metal2 s 376362 -960 376474 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 466 nsew signal input
flabel metal2 s 379674 -960 379786 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 467 nsew signal input
flabel metal2 s 382986 -960 383098 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 468 nsew signal input
flabel metal2 s 386298 -960 386410 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 469 nsew signal input
flabel metal2 s 389610 -960 389722 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 470 nsew signal input
flabel metal2 s 392922 -960 393034 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 471 nsew signal input
flabel metal2 s 396234 -960 396346 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 472 nsew signal input
flabel metal2 s 399546 -960 399658 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 473 nsew signal input
flabel metal2 s 402858 -960 402970 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 474 nsew signal input
flabel metal2 s 164394 -960 164506 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 475 nsew signal input
flabel metal2 s 406170 -960 406282 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 476 nsew signal input
flabel metal2 s 409482 -960 409594 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 477 nsew signal input
flabel metal2 s 412794 -960 412906 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 478 nsew signal input
flabel metal2 s 416106 -960 416218 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 479 nsew signal input
flabel metal2 s 419418 -960 419530 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 480 nsew signal input
flabel metal2 s 422730 -960 422842 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 481 nsew signal input
flabel metal2 s 426042 -960 426154 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 482 nsew signal input
flabel metal2 s 429354 -960 429466 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 483 nsew signal input
flabel metal2 s 432666 -960 432778 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 484 nsew signal input
flabel metal2 s 435978 -960 436090 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 485 nsew signal input
flabel metal2 s 167706 -960 167818 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 486 nsew signal input
flabel metal2 s 439290 -960 439402 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 487 nsew signal input
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 488 nsew signal input
flabel metal2 s 445914 -960 446026 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 489 nsew signal input
flabel metal2 s 449226 -960 449338 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 490 nsew signal input
flabel metal2 s 452538 -960 452650 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 491 nsew signal input
flabel metal2 s 455850 -960 455962 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 492 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 493 nsew signal input
flabel metal2 s 462474 -960 462586 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 494 nsew signal input
flabel metal2 s 465786 -960 465898 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 495 nsew signal input
flabel metal2 s 469098 -960 469210 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 496 nsew signal input
flabel metal2 s 171018 -960 171130 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 497 nsew signal input
flabel metal4 s -2316 -1244 -1696 705180 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -2316 -1244 586240 -624 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -2316 704560 586240 705180 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 585620 -1244 586240 705180 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 1794 -7964 2414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 37794 -7964 38414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 73794 -7964 74414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 109794 -7964 110414 98000 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 109794 152000 110414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 145794 -7964 146414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 181794 -7964 182414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 217794 -7964 218414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 253794 -7964 254414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 289794 -7964 290414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 325794 -7964 326414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 361794 -7964 362414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 397794 -7964 398414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 433794 -7964 434414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 469794 -7964 470414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 505794 -7964 506414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 541794 -7964 542414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s 577794 -7964 578414 711900 0 FreeSans 3840 90 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 2866 592960 3486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 38866 592960 39486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 74866 592960 75486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 110866 592960 111486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 146866 592960 147486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 182866 592960 183486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 218866 592960 219486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 254866 592960 255486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 290866 592960 291486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 326866 592960 327486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 362866 592960 363486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 398866 592960 399486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 434866 592960 435486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 470866 592960 471486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 506866 592960 507486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 542866 592960 543486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 578866 592960 579486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 614866 592960 615486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 650866 592960 651486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal5 s -9036 686866 592960 687486 0 FreeSans 2560 0 0 0 vccd1
port 498 nsew power bidirectional
flabel metal4 s -4236 -3164 -3616 707100 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -4236 -3164 588160 -2544 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -4236 706480 588160 707100 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 587540 -3164 588160 707100 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 10794 -7964 11414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 46794 -7964 47414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 82794 -7964 83414 98000 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 82794 152000 83414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 118794 -7964 119414 98000 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 118794 152000 119414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 154794 -7964 155414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 190794 -7964 191414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 226794 -7964 227414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 262794 -7964 263414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 298794 -7964 299414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 334794 -7964 335414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 370794 -7964 371414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 406794 -7964 407414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 442794 -7964 443414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 478794 -7964 479414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 514794 -7964 515414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s 550794 -7964 551414 711900 0 FreeSans 3840 90 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 11866 592960 12486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 47866 592960 48486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 83866 592960 84486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 119866 592960 120486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 155866 592960 156486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 191866 592960 192486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 227866 592960 228486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 263866 592960 264486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 299866 592960 300486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 335866 592960 336486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 371866 592960 372486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 407866 592960 408486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 443866 592960 444486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 479866 592960 480486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 515866 592960 516486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 551866 592960 552486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 587866 592960 588486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 623866 592960 624486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 659866 592960 660486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal5 s -9036 695866 592960 696486 0 FreeSans 2560 0 0 0 vccd2
port 499 nsew power bidirectional
flabel metal4 s -6156 -5084 -5536 709020 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -6156 -5084 590080 -4464 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -6156 708400 590080 709020 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 589460 -5084 590080 709020 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 19794 -7964 20414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 55794 -7964 56414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 91794 -7964 92414 98000 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 91794 152000 92414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 127794 -7964 128414 98000 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 127794 152000 128414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 163794 -7964 164414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 199794 -7964 200414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 235794 -7964 236414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 271794 -7964 272414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 307794 -7964 308414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 343794 -7964 344414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 379794 -7964 380414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 415794 -7964 416414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 451794 -7964 452414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 487794 -7964 488414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 523794 -7964 524414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s 559794 -7964 560414 711900 0 FreeSans 3840 90 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 20866 592960 21486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 56866 592960 57486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 92866 592960 93486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 128866 592960 129486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 164866 592960 165486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 200866 592960 201486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 236866 592960 237486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 272866 592960 273486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 308866 592960 309486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 344866 592960 345486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 380866 592960 381486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 416866 592960 417486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 452866 592960 453486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 488866 592960 489486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 524866 592960 525486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 560866 592960 561486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 596866 592960 597486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 632866 592960 633486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal5 s -9036 668866 592960 669486 0 FreeSans 2560 0 0 0 vdda1
port 500 nsew power bidirectional
flabel metal4 s -8076 -7004 -7456 710940 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -8076 -7004 592000 -6384 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -8076 710320 592000 710940 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 591380 -7004 592000 710940 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 28794 -7964 29414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 64794 -7964 65414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 100794 -7964 101414 98000 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 100794 152000 101414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 136794 -7964 137414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 172794 -7964 173414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 208794 -7964 209414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 244794 -7964 245414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 280794 -7964 281414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 316794 -7964 317414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 352794 -7964 353414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 388794 -7964 389414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 424794 -7964 425414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 460794 -7964 461414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 496794 -7964 497414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 532794 -7964 533414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s 568794 -7964 569414 711900 0 FreeSans 3840 90 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 29866 592960 30486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 65866 592960 66486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 101866 592960 102486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 137866 592960 138486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 173866 592960 174486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 209866 592960 210486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 245866 592960 246486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 281866 592960 282486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 317866 592960 318486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 353866 592960 354486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 389866 592960 390486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 425866 592960 426486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 461866 592960 462486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 497866 592960 498486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 533866 592960 534486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 569866 592960 570486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 605866 592960 606486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 641866 592960 642486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal5 s -9036 677866 592960 678486 0 FreeSans 2560 0 0 0 vdda2
port 501 nsew power bidirectional
flabel metal4 s -7116 -6044 -6496 709980 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -7116 -6044 591040 -5424 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -7116 709360 591040 709980 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 590420 -6044 591040 709980 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 24294 -7964 24914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 60294 -7964 60914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 96294 -7964 96914 98000 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 96294 152000 96914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 132294 -7964 132914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 168294 -7964 168914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 204294 -7964 204914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 240294 -7964 240914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 276294 -7964 276914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 312294 -7964 312914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 348294 -7964 348914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 384294 -7964 384914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 420294 -7964 420914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 456294 -7964 456914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 492294 -7964 492914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 528294 -7964 528914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s 564294 -7964 564914 711900 0 FreeSans 3840 90 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 25366 592960 25986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 61366 592960 61986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 97366 592960 97986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 133366 592960 133986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 169366 592960 169986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 205366 592960 205986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 241366 592960 241986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 277366 592960 277986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 313366 592960 313986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 349366 592960 349986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 385366 592960 385986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 421366 592960 421986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 457366 592960 457986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 493366 592960 493986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 529366 592960 529986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 565366 592960 565986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 601366 592960 601986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 637366 592960 637986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal5 s -9036 673366 592960 673986 0 FreeSans 2560 0 0 0 vssa1
port 502 nsew ground bidirectional
flabel metal4 s -9036 -7964 -8416 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 -7964 592960 -7344 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 711280 592960 711900 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 592340 -7964 592960 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 33294 -7964 33914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 69294 -7964 69914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 105294 -7964 105914 98000 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 105294 152000 105914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 141294 -7964 141914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 177294 -7964 177914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 213294 -7964 213914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 249294 -7964 249914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 285294 -7964 285914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 321294 -7964 321914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 357294 -7964 357914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 393294 -7964 393914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 429294 -7964 429914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 465294 -7964 465914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 501294 -7964 501914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 537294 -7964 537914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s 573294 -7964 573914 711900 0 FreeSans 3840 90 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 34366 592960 34986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 70366 592960 70986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 106366 592960 106986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 142366 592960 142986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 178366 592960 178986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 214366 592960 214986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 250366 592960 250986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 286366 592960 286986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 322366 592960 322986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 358366 592960 358986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 394366 592960 394986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 430366 592960 430986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 466366 592960 466986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 502366 592960 502986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 538366 592960 538986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 574366 592960 574986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 610366 592960 610986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 646366 592960 646986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal5 s -9036 682366 592960 682986 0 FreeSans 2560 0 0 0 vssa2
port 503 nsew ground bidirectional
flabel metal4 s -3276 -2204 -2656 706140 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -3276 -2204 587200 -1584 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -3276 705520 587200 706140 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 586580 -2204 587200 706140 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 6294 -7964 6914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 42294 -7964 42914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 78294 -7964 78914 98000 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 78294 152000 78914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 114294 -7964 114914 98000 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 114294 152000 114914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 150294 -7964 150914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 186294 -7964 186914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 222294 -7964 222914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 258294 -7964 258914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 294294 -7964 294914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 330294 -7964 330914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 366294 -7964 366914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 402294 -7964 402914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 438294 -7964 438914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 474294 -7964 474914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 510294 -7964 510914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 546294 -7964 546914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s 582294 -7964 582914 711900 0 FreeSans 3840 90 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 7366 592960 7986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 43366 592960 43986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 79366 592960 79986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 115366 592960 115986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 151366 592960 151986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 187366 592960 187986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 223366 592960 223986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 259366 592960 259986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 295366 592960 295986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 331366 592960 331986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 367366 592960 367986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 403366 592960 403986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 439366 592960 439986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 475366 592960 475986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 511366 592960 511986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 547366 592960 547986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 583366 592960 583986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 619366 592960 619986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 655366 592960 655986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal5 s -9036 691366 592960 691986 0 FreeSans 2560 0 0 0 vssd1
port 504 nsew ground bidirectional
flabel metal4 s -5196 -4124 -4576 708060 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -5196 -4124 589120 -3504 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -5196 707440 589120 708060 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 588500 -4124 589120 708060 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 15294 -7964 15914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 51294 -7964 51914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 87294 -7964 87914 98000 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 87294 152000 87914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 123294 -7964 123914 98000 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 123294 152000 123914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 159294 -7964 159914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 195294 -7964 195914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 231294 -7964 231914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 267294 -7964 267914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 303294 -7964 303914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 339294 -7964 339914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 375294 -7964 375914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 411294 -7964 411914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 447294 -7964 447914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 483294 -7964 483914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 519294 -7964 519914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal4 s 555294 -7964 555914 711900 0 FreeSans 3840 90 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 16366 592960 16986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 52366 592960 52986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 88366 592960 88986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 124366 592960 124986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 160366 592960 160986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 196366 592960 196986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 232366 592960 232986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 268366 592960 268986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 304366 592960 304986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 340366 592960 340986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 376366 592960 376986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 412366 592960 412986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 448366 592960 448986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 484366 592960 484986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 520366 592960 520986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 556366 592960 556986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 592366 592960 592986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 628366 592960 628986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 664366 592960 664986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal5 s -9036 700366 592960 700986 0 FreeSans 2560 0 0 0 vssd2
port 505 nsew ground bidirectional
flabel metal2 s 21978 -960 22090 480 0 FreeSans 448 90 0 0 wb_clk_i
port 506 nsew signal input
flabel metal2 s 23082 -960 23194 480 0 FreeSans 448 90 0 0 wb_rst_i
port 507 nsew signal input
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 508 nsew signal tristate
flabel metal2 s 28602 -960 28714 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 509 nsew signal input
flabel metal2 s 66138 -960 66250 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 510 nsew signal input
flabel metal2 s 69450 -960 69562 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 511 nsew signal input
flabel metal2 s 72762 -960 72874 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 512 nsew signal input
flabel metal2 s 76074 -960 76186 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 513 nsew signal input
flabel metal2 s 79386 -960 79498 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 514 nsew signal input
flabel metal2 s 82698 -960 82810 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 515 nsew signal input
flabel metal2 s 86010 -960 86122 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 516 nsew signal input
flabel metal2 s 89322 -960 89434 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 517 nsew signal input
flabel metal2 s 92634 -960 92746 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 518 nsew signal input
flabel metal2 s 95946 -960 96058 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 519 nsew signal input
flabel metal2 s 33018 -960 33130 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 520 nsew signal input
flabel metal2 s 99258 -960 99370 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 521 nsew signal input
flabel metal2 s 102570 -960 102682 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 522 nsew signal input
flabel metal2 s 105882 -960 105994 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 523 nsew signal input
flabel metal2 s 109194 -960 109306 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 524 nsew signal input
flabel metal2 s 112506 -960 112618 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 525 nsew signal input
flabel metal2 s 115818 -960 115930 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 526 nsew signal input
flabel metal2 s 119130 -960 119242 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 527 nsew signal input
flabel metal2 s 122442 -960 122554 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 528 nsew signal input
flabel metal2 s 125754 -960 125866 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 529 nsew signal input
flabel metal2 s 129066 -960 129178 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 530 nsew signal input
flabel metal2 s 37434 -960 37546 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 531 nsew signal input
flabel metal2 s 132378 -960 132490 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 532 nsew signal input
flabel metal2 s 135690 -960 135802 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 533 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 534 nsew signal input
flabel metal2 s 46266 -960 46378 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 535 nsew signal input
flabel metal2 s 49578 -960 49690 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 536 nsew signal input
flabel metal2 s 52890 -960 53002 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 537 nsew signal input
flabel metal2 s 56202 -960 56314 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 538 nsew signal input
flabel metal2 s 59514 -960 59626 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 539 nsew signal input
flabel metal2 s 62826 -960 62938 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 540 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 541 nsew signal input
flabel metal2 s 29706 -960 29818 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 542 nsew signal input
flabel metal2 s 67242 -960 67354 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 543 nsew signal input
flabel metal2 s 70554 -960 70666 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 544 nsew signal input
flabel metal2 s 73866 -960 73978 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 545 nsew signal input
flabel metal2 s 77178 -960 77290 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 546 nsew signal input
flabel metal2 s 80490 -960 80602 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 547 nsew signal input
flabel metal2 s 83802 -960 83914 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 548 nsew signal input
flabel metal2 s 87114 -960 87226 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 549 nsew signal input
flabel metal2 s 90426 -960 90538 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 550 nsew signal input
flabel metal2 s 93738 -960 93850 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 551 nsew signal input
flabel metal2 s 97050 -960 97162 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 552 nsew signal input
flabel metal2 s 34122 -960 34234 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 553 nsew signal input
flabel metal2 s 100362 -960 100474 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 554 nsew signal input
flabel metal2 s 103674 -960 103786 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 555 nsew signal input
flabel metal2 s 106986 -960 107098 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 556 nsew signal input
flabel metal2 s 110298 -960 110410 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 557 nsew signal input
flabel metal2 s 113610 -960 113722 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 558 nsew signal input
flabel metal2 s 116922 -960 117034 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 559 nsew signal input
flabel metal2 s 120234 -960 120346 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 560 nsew signal input
flabel metal2 s 123546 -960 123658 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 561 nsew signal input
flabel metal2 s 126858 -960 126970 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 562 nsew signal input
flabel metal2 s 130170 -960 130282 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 563 nsew signal input
flabel metal2 s 38538 -960 38650 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 564 nsew signal input
flabel metal2 s 133482 -960 133594 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 565 nsew signal input
flabel metal2 s 136794 -960 136906 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 566 nsew signal input
flabel metal2 s 42954 -960 43066 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 567 nsew signal input
flabel metal2 s 47370 -960 47482 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 568 nsew signal input
flabel metal2 s 50682 -960 50794 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 569 nsew signal input
flabel metal2 s 53994 -960 54106 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 570 nsew signal input
flabel metal2 s 57306 -960 57418 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 571 nsew signal input
flabel metal2 s 60618 -960 60730 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 572 nsew signal input
flabel metal2 s 63930 -960 64042 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 573 nsew signal input
flabel metal2 s 30810 -960 30922 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 574 nsew signal tristate
flabel metal2 s 68346 -960 68458 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 575 nsew signal tristate
flabel metal2 s 71658 -960 71770 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 576 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 577 nsew signal tristate
flabel metal2 s 78282 -960 78394 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 578 nsew signal tristate
flabel metal2 s 81594 -960 81706 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 579 nsew signal tristate
flabel metal2 s 84906 -960 85018 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 580 nsew signal tristate
flabel metal2 s 88218 -960 88330 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 581 nsew signal tristate
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 582 nsew signal tristate
flabel metal2 s 94842 -960 94954 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 583 nsew signal tristate
flabel metal2 s 98154 -960 98266 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 584 nsew signal tristate
flabel metal2 s 35226 -960 35338 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 585 nsew signal tristate
flabel metal2 s 101466 -960 101578 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 586 nsew signal tristate
flabel metal2 s 104778 -960 104890 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 587 nsew signal tristate
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 588 nsew signal tristate
flabel metal2 s 111402 -960 111514 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 589 nsew signal tristate
flabel metal2 s 114714 -960 114826 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 590 nsew signal tristate
flabel metal2 s 118026 -960 118138 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 591 nsew signal tristate
flabel metal2 s 121338 -960 121450 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 592 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 593 nsew signal tristate
flabel metal2 s 127962 -960 128074 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 594 nsew signal tristate
flabel metal2 s 131274 -960 131386 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 595 nsew signal tristate
flabel metal2 s 39642 -960 39754 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 596 nsew signal tristate
flabel metal2 s 134586 -960 134698 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 597 nsew signal tristate
flabel metal2 s 137898 -960 138010 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 598 nsew signal tristate
flabel metal2 s 44058 -960 44170 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 599 nsew signal tristate
flabel metal2 s 48474 -960 48586 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 600 nsew signal tristate
flabel metal2 s 51786 -960 51898 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 601 nsew signal tristate
flabel metal2 s 55098 -960 55210 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 602 nsew signal tristate
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 603 nsew signal tristate
flabel metal2 s 61722 -960 61834 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 604 nsew signal tristate
flabel metal2 s 65034 -960 65146 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 605 nsew signal tristate
flabel metal2 s 31914 -960 32026 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 606 nsew signal input
flabel metal2 s 36330 -960 36442 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 607 nsew signal input
flabel metal2 s 40746 -960 40858 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 608 nsew signal input
flabel metal2 s 45162 -960 45274 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 609 nsew signal input
flabel metal2 s 26394 -960 26506 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 610 nsew signal input
flabel metal2 s 27498 -960 27610 480 0 FreeSans 448 90 0 0 wbs_we_i
port 611 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
